magic
tech sky130A
magscale 1 2
timestamp 1771143426
<< nwell >>
rect -4000 -10000 9200 -8700
rect -4000 -11200 900 -10000
rect -4000 -12900 -2200 -11200
rect 4300 -11200 9200 -10000
rect -4000 -14460 700 -12900
rect 7400 -12900 9200 -11200
rect 4500 -14460 9200 -12900
rect -4000 -14700 9200 -14460
<< pwell >>
rect 1000 -11300 4200 -10100
rect -2100 -12800 7300 -11300
rect 800 -14400 4400 -12800
<< psubdiff >>
rect 1000 -10120 4200 -10100
rect 1000 -10180 1120 -10120
rect 4100 -10180 4200 -10120
rect 1000 -10200 4200 -10180
rect 1000 -10220 1100 -10200
rect 1000 -11280 1020 -10220
rect 1080 -11280 1100 -10220
rect 1000 -11300 1100 -11280
rect -2100 -11320 1100 -11300
rect -2100 -11380 -1980 -11320
rect 980 -11380 1100 -11320
rect -2100 -11400 1100 -11380
rect 4100 -10220 4200 -10200
rect 4100 -11280 4120 -10220
rect 4180 -11280 4200 -10220
rect 4100 -11300 4200 -11280
rect 4100 -11320 7300 -11300
rect 4100 -11380 4220 -11320
rect 7180 -11380 7300 -11320
rect 4100 -11400 7300 -11380
rect -2100 -11420 -2000 -11400
rect -2100 -12680 -2080 -11420
rect -2020 -12680 -2000 -11420
rect -2100 -12700 -2000 -12680
rect 7200 -11420 7300 -11400
rect 7200 -12680 7220 -11420
rect 7280 -12680 7300 -11420
rect 7200 -12700 7300 -12680
rect -2100 -12720 900 -12700
rect -2100 -12780 -1980 -12720
rect 780 -12780 900 -12720
rect -2100 -12800 900 -12780
rect 800 -12820 900 -12800
rect 800 -14280 820 -12820
rect 880 -14280 900 -12820
rect 800 -14300 900 -14280
rect 4300 -12720 7300 -12700
rect 4300 -12780 4420 -12720
rect 7180 -12780 7300 -12720
rect 4300 -12800 7300 -12780
rect 4300 -12820 4400 -12800
rect 4300 -14280 4320 -12820
rect 4380 -14280 4400 -12820
rect 4300 -14300 4400 -14280
rect 800 -14320 4400 -14300
rect 800 -14380 900 -14320
rect 4280 -14380 4400 -14320
rect 800 -14400 4400 -14380
<< nsubdiff >>
rect -3900 -8820 9100 -8800
rect -3900 -8880 -3780 -8820
rect 8980 -8880 9100 -8820
rect -3900 -8900 9100 -8880
rect -3900 -8920 -3800 -8900
rect -3900 -14480 -3880 -8920
rect -3820 -14480 -3800 -8920
rect 9000 -8940 9100 -8900
rect -3900 -14500 -3800 -14480
rect 9000 -14500 9020 -8940
rect 9080 -14500 9100 -8940
rect -3900 -14520 9100 -14500
rect -3900 -14580 -3780 -14520
rect 8980 -14580 9100 -14520
rect -3900 -14600 9100 -14580
<< psubdiffcont >>
rect 1120 -10180 4100 -10120
rect 1020 -11280 1080 -10220
rect -1980 -11380 980 -11320
rect 4120 -11280 4180 -10220
rect 4220 -11380 7180 -11320
rect -2080 -12680 -2020 -11420
rect 7220 -12680 7280 -11420
rect -1980 -12780 780 -12720
rect 820 -14280 880 -12820
rect 4420 -12780 7180 -12720
rect 4320 -14280 4380 -12820
rect 900 -14380 4280 -14320
<< nsubdiffcont >>
rect -3780 -8880 8980 -8820
rect -3880 -14480 -3820 -8920
rect 9020 -14500 9080 -8940
rect -3780 -14580 8980 -14520
<< locali >>
rect -3900 -8820 9100 -8800
rect -3900 -8880 -3780 -8820
rect 8980 -8880 9100 -8820
rect -3900 -8900 9100 -8880
rect -3900 -8920 2540 -8900
rect -3900 -14480 -3880 -8920
rect -3820 -8980 2540 -8920
rect 2620 -8940 9100 -8900
rect 2620 -8980 9020 -8940
rect -3820 -9100 9020 -8980
rect -3820 -9940 -1800 -9100
rect -1500 -9880 -1360 -9100
rect -880 -9880 -740 -9100
rect -260 -9880 -120 -9100
rect 360 -9880 500 -9100
rect 840 -9140 4340 -9100
rect 840 -9900 1060 -9140
rect 1420 -9780 1520 -9140
rect 2040 -9780 2140 -9140
rect 2520 -9900 2660 -9140
rect 3020 -9780 3120 -9140
rect 3640 -9780 3740 -9140
rect 4120 -9900 4340 -9140
rect 4700 -9860 4840 -9100
rect 5320 -9860 5460 -9100
rect 5940 -9860 6080 -9100
rect 6560 -9860 6700 -9100
rect -3820 -10020 -3100 -9940
rect -3020 -10020 -1800 -9940
rect -3820 -10040 -1800 -10020
rect 800 -10000 4400 -9900
rect 800 -10040 900 -10000
rect -3820 -10200 900 -10040
rect 4300 -10060 4400 -10000
rect 7000 -10060 9020 -9100
rect -3820 -11100 -3640 -10200
rect -960 -10340 900 -10200
rect -3300 -11100 -3160 -10380
rect -2680 -11100 -2540 -10380
rect -2060 -11100 -1920 -10380
rect -1440 -11100 -1300 -10380
rect -940 -11100 -660 -10340
rect -300 -10980 -160 -10340
rect 320 -10980 460 -10340
rect 800 -11100 900 -10340
rect -3820 -11200 900 -11100
rect 1000 -10120 4200 -10100
rect 1000 -10180 1120 -10120
rect 4100 -10180 4200 -10120
rect 1000 -10220 4200 -10180
rect -3820 -12900 -2180 -11200
rect 1000 -11280 1020 -10220
rect 1080 -10440 4120 -10220
rect 1080 -10940 2240 -10440
rect 2960 -10940 4120 -10440
rect 1080 -11220 4120 -10940
rect 1080 -11280 2180 -11220
rect 1000 -11300 2180 -11280
rect -2100 -11320 2180 -11300
rect -2100 -11380 -1980 -11320
rect 980 -11380 2180 -11320
rect -2100 -11420 2180 -11380
rect -2100 -12680 -2080 -11420
rect -2020 -11540 2180 -11420
rect -2020 -12440 -1740 -11540
rect -900 -11620 2180 -11540
rect -1380 -12440 -1260 -11820
rect -900 -12440 -660 -11620
rect -300 -12380 -180 -11620
rect -120 -12160 2180 -11620
rect 2546 -11994 2636 -11220
rect 3020 -11280 4120 -11220
rect 4180 -11280 4200 -10220
rect 4300 -10200 9020 -10060
rect 4300 -10340 6140 -10200
rect 4300 -11100 4400 -10340
rect 4700 -10980 4840 -10340
rect 5340 -10980 5480 -10340
rect 5820 -11100 6140 -10340
rect 6500 -11100 6640 -10380
rect 7120 -11100 7260 -10380
rect 7740 -11100 7880 -10380
rect 8360 -11100 8500 -10380
rect 8840 -11100 9020 -10200
rect 4300 -11200 9020 -11100
rect 3020 -11300 4200 -11280
rect 3020 -11320 7300 -11300
rect 3020 -11380 4220 -11320
rect 7180 -11380 7300 -11320
rect 3020 -11420 7300 -11380
rect 3020 -11494 7220 -11420
rect 3020 -11540 4768 -11494
rect 3020 -11940 4760 -11540
rect 5080 -11584 7220 -11494
rect 5080 -11620 6060 -11584
rect 5080 -11940 5240 -11620
rect 3020 -12160 5240 -11940
rect -120 -12340 5240 -12160
rect -2020 -12560 -660 -12440
rect -120 -12540 1140 -12340
rect -260 -12560 1140 -12540
rect -2020 -12680 1140 -12560
rect -2100 -12720 1140 -12680
rect -2100 -12780 -1980 -12720
rect 780 -12780 1140 -12720
rect -2100 -12800 1140 -12780
rect 800 -12820 1140 -12800
rect -3820 -14460 700 -12900
rect 800 -14280 820 -12820
rect 880 -13620 1140 -12820
rect 880 -13680 900 -13620
rect 960 -13680 1140 -13620
rect 880 -13740 1140 -13680
rect 880 -13800 900 -13740
rect 960 -13800 1140 -13740
rect 880 -14040 1140 -13800
rect 1660 -14040 1760 -12340
rect 2260 -14040 2360 -12340
rect 2860 -14040 2960 -12340
rect 3460 -14040 3560 -12340
rect 4060 -12540 5240 -12340
rect 5780 -12440 6060 -11620
rect 6420 -12440 6540 -11820
rect 6900 -12440 7220 -11584
rect 5780 -12540 7220 -12440
rect 4060 -12680 7220 -12540
rect 7280 -12680 7300 -11420
rect 4060 -12720 7300 -12680
rect 4060 -12780 4420 -12720
rect 7180 -12780 7300 -12720
rect 4060 -12800 7300 -12780
rect 4060 -12820 4400 -12800
rect 4060 -14040 4320 -12820
rect 880 -14140 4320 -14040
rect 880 -14200 900 -14140
rect 960 -14200 4320 -14140
rect 880 -14240 4320 -14200
rect 880 -14280 900 -14240
rect 800 -14300 900 -14280
rect 960 -14300 4240 -14240
rect 4300 -14280 4320 -14240
rect 4380 -14280 4400 -12820
rect 7400 -12900 9020 -11200
rect 4300 -14300 4400 -14280
rect 800 -14320 4400 -14300
rect 800 -14380 900 -14320
rect 4280 -14380 4400 -14320
rect 800 -14400 4400 -14380
rect 4500 -14460 9020 -12900
rect -3820 -14480 9020 -14460
rect -3900 -14500 9020 -14480
rect 9080 -14500 9100 -8940
rect -3900 -14520 9100 -14500
rect -3900 -14580 -3780 -14520
rect 8980 -14580 9100 -14520
rect -3900 -14600 9100 -14580
<< viali >>
rect -3100 -10020 -3020 -9940
rect 900 -13680 960 -13620
rect 900 -13800 960 -13740
rect 900 -14200 960 -14140
rect 900 -14300 960 -14240
rect 4240 -14300 4300 -14240
<< metal1 >>
rect 2480 -8480 2680 -8460
rect 2480 -8560 2540 -8480
rect 2620 -8560 2680 -8480
rect 2480 -8580 2680 -8560
rect 2480 -8660 2540 -8580
rect 2620 -8660 2680 -8580
rect 2500 -8700 2660 -8660
rect 2500 -8780 2540 -8700
rect 2620 -8780 2660 -8700
rect 2500 -8800 2660 -8780
rect 2500 -8880 2540 -8800
rect 2620 -8880 2660 -8800
rect 2500 -8900 2660 -8880
rect 2500 -8980 2540 -8900
rect 2620 -8980 2660 -8900
rect 2500 -9000 2660 -8980
rect 2500 -9080 2540 -9000
rect 2620 -9080 2660 -9000
rect 2500 -9100 2660 -9080
rect 2500 -9180 2540 -9100
rect 2620 -9180 2660 -9100
rect 2500 -9200 2660 -9180
rect -1800 -9420 -1680 -9400
rect -1800 -9500 -1780 -9420
rect -1700 -9500 -1680 -9420
rect -1800 -9560 -1680 -9500
rect -3400 -9934 -3000 -9600
rect -1800 -9640 -1780 -9560
rect -1700 -9640 -1680 -9560
rect -1800 -9660 -1680 -9640
rect -1180 -9420 -1060 -9400
rect -1180 -9500 -1160 -9420
rect -1080 -9500 -1060 -9420
rect -1180 -9560 -1060 -9500
rect -1180 -9640 -1160 -9560
rect -1080 -9640 -1060 -9560
rect -1180 -9660 -1060 -9640
rect -560 -9420 -440 -9400
rect -560 -9500 -540 -9420
rect -460 -9500 -440 -9420
rect -560 -9560 -440 -9500
rect -560 -9640 -540 -9560
rect -460 -9640 -440 -9560
rect -560 -9660 -440 -9640
rect 40 -9420 160 -9400
rect 40 -9500 60 -9420
rect 140 -9500 160 -9420
rect 40 -9560 160 -9500
rect 40 -9640 60 -9560
rect 140 -9640 160 -9560
rect 40 -9660 160 -9640
rect 640 -9420 760 -9400
rect 640 -9500 660 -9420
rect 740 -9500 760 -9420
rect 640 -9560 760 -9500
rect 640 -9640 660 -9560
rect 740 -9640 760 -9560
rect 640 -9660 760 -9640
rect 1140 -9820 1240 -9240
rect 1740 -9440 1840 -9240
rect 1740 -9480 1860 -9440
rect 1740 -9540 1780 -9480
rect 1840 -9540 1860 -9480
rect 1740 -9580 1860 -9540
rect 2340 -9480 2440 -9240
rect 2500 -9280 2540 -9200
rect 2620 -9280 2660 -9200
rect 2500 -9300 2660 -9280
rect 2500 -9380 2540 -9300
rect 2620 -9380 2660 -9300
rect 2500 -9400 2660 -9380
rect 4440 -9420 4560 -9400
rect 2340 -9540 2360 -9480
rect 2420 -9540 2440 -9480
rect 1740 -9820 1840 -9580
rect 2340 -9820 2440 -9540
rect 2720 -9480 2820 -9440
rect 2720 -9540 2740 -9480
rect 2800 -9540 2820 -9480
rect 2720 -9580 2820 -9540
rect 3320 -9480 3420 -9440
rect 3320 -9540 3340 -9480
rect 3400 -9540 3420 -9480
rect 3320 -9580 3420 -9540
rect 3940 -9480 4040 -9440
rect 3940 -9540 3960 -9480
rect 4020 -9540 4040 -9480
rect 3940 -9580 4040 -9540
rect 4440 -9500 4460 -9420
rect 4540 -9500 4560 -9420
rect 4440 -9560 4560 -9500
rect 4440 -9640 4460 -9560
rect 4540 -9640 4560 -9560
rect 4440 -9660 4560 -9640
rect 5020 -9420 5140 -9400
rect 5020 -9500 5040 -9420
rect 5120 -9500 5140 -9420
rect 5020 -9560 5140 -9500
rect 5020 -9640 5040 -9560
rect 5120 -9640 5140 -9560
rect 5020 -9660 5140 -9640
rect 5640 -9420 5760 -9400
rect 5640 -9500 5660 -9420
rect 5740 -9500 5760 -9420
rect 5640 -9560 5760 -9500
rect 5640 -9640 5660 -9560
rect 5740 -9640 5760 -9560
rect 5640 -9660 5760 -9640
rect 6260 -9420 6380 -9400
rect 6260 -9500 6280 -9420
rect 6360 -9500 6380 -9420
rect 6260 -9560 6380 -9500
rect 6260 -9640 6280 -9560
rect 6360 -9640 6380 -9560
rect 6260 -9660 6380 -9640
rect 6860 -9420 6980 -9400
rect 6860 -9500 6880 -9420
rect 6960 -9500 6980 -9420
rect 6860 -9560 6980 -9500
rect 6860 -9640 6880 -9560
rect 6960 -9640 6980 -9560
rect 6860 -9660 6980 -9640
rect 1140 -9900 4000 -9820
rect 8200 -9934 8600 -9600
rect -3520 -9940 -960 -9934
rect -760 -9940 2500 -9934
rect 2580 -9940 2620 -9934
rect 2700 -9940 5900 -9934
rect 6100 -9940 8710 -9934
rect -3520 -10020 -3380 -9940
rect -3300 -10020 -3100 -9940
rect -3020 -10000 3300 -9940
rect 3360 -10000 8220 -9940
rect -3020 -10020 8220 -10000
rect 8300 -10020 8500 -9940
rect 8580 -10020 8710 -9940
rect -3520 -10080 3300 -10020
rect 3360 -10080 8710 -10020
rect -3520 -10100 8710 -10080
rect -3520 -10180 -3380 -10100
rect -3300 -10180 -3100 -10100
rect -3020 -10160 8220 -10100
rect -3020 -10180 3300 -10160
rect -3520 -10220 3300 -10180
rect 3360 -10180 8220 -10160
rect 8300 -10180 8500 -10100
rect 8580 -10180 8710 -10100
rect 3360 -10220 8710 -10180
rect -3520 -10240 8710 -10220
rect -3520 -10300 3300 -10240
rect 3360 -10300 8710 -10240
rect -3520 -10316 8710 -10300
rect -1120 -10320 -620 -10316
rect 2500 -10320 2700 -10316
rect 5760 -10320 6220 -10316
rect 2120 -10380 2460 -10360
rect 1760 -10420 1860 -10380
rect -600 -10460 -460 -10440
rect -600 -10560 -580 -10460
rect -480 -10560 -460 -10460
rect -3560 -10600 -3440 -10580
rect -3560 -10680 -3540 -10600
rect -3460 -10680 -3440 -10600
rect -3560 -10740 -3440 -10680
rect -3560 -10820 -3540 -10740
rect -3460 -10820 -3440 -10740
rect -3560 -10840 -3440 -10820
rect -2980 -10600 -2860 -10580
rect -2980 -10680 -2960 -10600
rect -2880 -10680 -2860 -10600
rect -2980 -10740 -2860 -10680
rect -2980 -10820 -2960 -10740
rect -2880 -10820 -2860 -10740
rect -2980 -10840 -2860 -10820
rect -2360 -10600 -2240 -10580
rect -2360 -10680 -2340 -10600
rect -2260 -10680 -2240 -10600
rect -2360 -10740 -2240 -10680
rect -2360 -10820 -2340 -10740
rect -2260 -10820 -2240 -10740
rect -2360 -10840 -2240 -10820
rect -1740 -10600 -1620 -10580
rect -1740 -10680 -1720 -10600
rect -1640 -10680 -1620 -10600
rect -1740 -10740 -1620 -10680
rect -1740 -10820 -1720 -10740
rect -1640 -10820 -1620 -10740
rect -1740 -10840 -1620 -10820
rect -1160 -10600 -1040 -10580
rect -1160 -10680 -1140 -10600
rect -1060 -10680 -1040 -10600
rect -1160 -10740 -1040 -10680
rect -1160 -10820 -1140 -10740
rect -1060 -10820 -1040 -10740
rect -1160 -10840 -1040 -10820
rect -600 -10660 -460 -10560
rect -600 -10760 -580 -10660
rect -480 -10760 -460 -10660
rect -600 -10860 -460 -10760
rect -600 -10960 -580 -10860
rect -480 -10960 -460 -10860
rect -600 -10980 -460 -10960
rect 20 -10660 160 -10440
rect 20 -10760 40 -10660
rect 140 -10760 160 -10660
rect 20 -10980 160 -10760
rect 620 -10660 760 -10440
rect 620 -10760 640 -10660
rect 740 -10760 760 -10660
rect 620 -10980 760 -10760
rect 1760 -10480 1780 -10420
rect 1840 -10480 1860 -10420
rect 2120 -10440 2140 -10380
rect 2200 -10440 2240 -10380
rect 2300 -10440 2380 -10380
rect 2440 -10440 2460 -10380
rect 2120 -10460 2460 -10440
rect 1760 -10780 1860 -10480
rect 2380 -10560 2460 -10460
rect 2500 -10380 2700 -10360
rect 2500 -10440 2520 -10380
rect 2580 -10440 2620 -10380
rect 2680 -10440 2700 -10380
rect 2500 -10480 2700 -10440
rect 2500 -10540 2520 -10480
rect 2580 -10540 2620 -10480
rect 2680 -10540 2700 -10480
rect 2500 -10560 2700 -10540
rect 2740 -10380 3080 -10360
rect 2740 -10440 2760 -10380
rect 2820 -10440 2900 -10380
rect 2960 -10440 3000 -10380
rect 3060 -10440 3080 -10380
rect 2740 -10460 3080 -10440
rect 2740 -10560 2820 -10460
rect 1760 -10840 1780 -10780
rect 1840 -10840 1860 -10780
rect 1760 -10860 1860 -10840
rect 2320 -10780 2400 -10760
rect 2320 -10840 2340 -10780
rect 2320 -10860 2400 -10840
rect 2440 -10900 2540 -10600
rect 2580 -10620 2640 -10600
rect 2580 -10700 2640 -10680
rect 2680 -10900 2780 -10600
rect 2820 -10780 2900 -10760
rect 2880 -10840 2900 -10780
rect 2820 -10860 2900 -10840
rect 1760 -10940 3380 -10900
rect 1760 -11000 1800 -10940
rect 1860 -11000 3280 -10940
rect 3340 -11000 3380 -10940
rect 4400 -11032 4520 -10440
rect 5020 -11032 5140 -10440
rect 5640 -11032 5760 -10440
rect 6220 -10600 6340 -10580
rect 6220 -10680 6240 -10600
rect 6320 -10680 6340 -10600
rect 6220 -10740 6340 -10680
rect 6220 -10820 6240 -10740
rect 6320 -10820 6340 -10740
rect 6220 -10840 6340 -10820
rect 6820 -10600 6940 -10580
rect 6820 -10680 6840 -10600
rect 6920 -10680 6940 -10600
rect 6820 -10740 6940 -10680
rect 6820 -10820 6840 -10740
rect 6920 -10820 6940 -10740
rect 6820 -10840 6940 -10820
rect 7440 -10600 7560 -10580
rect 7440 -10680 7460 -10600
rect 7540 -10680 7560 -10600
rect 7440 -10740 7560 -10680
rect 7440 -10820 7460 -10740
rect 7540 -10820 7560 -10740
rect 7440 -10840 7560 -10820
rect 8060 -10600 8180 -10580
rect 8060 -10680 8080 -10600
rect 8160 -10680 8180 -10600
rect 8060 -10740 8180 -10680
rect 8060 -10820 8080 -10740
rect 8160 -10820 8180 -10740
rect 8060 -10840 8180 -10820
rect 8620 -10600 8740 -10580
rect 8620 -10680 8640 -10600
rect 8720 -10680 8740 -10600
rect 8620 -10740 8740 -10680
rect 8620 -10820 8640 -10740
rect 8720 -10820 8740 -10740
rect 8620 -10840 8740 -10820
rect -500 -11040 20 -11032
rect 140 -11040 640 -11032
rect 760 -11040 5844 -11032
rect -500 -11246 5844 -11040
rect 200 -11300 280 -11246
rect -1640 -11660 -960 -11300
rect 20 -11340 280 -11300
rect 2320 -11320 2880 -11246
rect 20 -11400 40 -11340
rect 100 -11400 200 -11340
rect 260 -11400 280 -11340
rect 20 -11440 280 -11400
rect 4952 -11540 5034 -11246
rect 2240 -11600 2340 -11580
rect 2240 -11660 2260 -11600
rect 2320 -11660 2340 -11600
rect -1620 -11700 -1040 -11660
rect 2240 -11700 2340 -11660
rect -600 -11740 -460 -11720
rect -600 -11840 -580 -11740
rect -480 -11840 -460 -11740
rect 2240 -11760 2260 -11700
rect 2320 -11760 2340 -11700
rect 2240 -11780 2340 -11760
rect 2860 -11600 2960 -11580
rect 2860 -11660 2880 -11600
rect 2940 -11660 2960 -11600
rect 2860 -11700 2960 -11660
rect 2860 -11760 2880 -11700
rect 2940 -11760 2960 -11700
rect 2860 -11780 2960 -11760
rect -600 -11880 -460 -11840
rect -1700 -11940 -1580 -11920
rect -2600 -12020 -2200 -12000
rect -2600 -12100 -2580 -12020
rect -2500 -12100 -2300 -12020
rect -2220 -12100 -2200 -12020
rect -2600 -12500 -2200 -12100
rect -1700 -12020 -1680 -11940
rect -1600 -12020 -1580 -11940
rect -1700 -12080 -1580 -12020
rect -1700 -12160 -1680 -12080
rect -1600 -12160 -1580 -12080
rect -1700 -12180 -1580 -12160
rect -1100 -11940 -980 -11920
rect -1100 -12020 -1080 -11940
rect -1000 -12020 -980 -11940
rect -1100 -12080 -980 -12020
rect -1100 -12160 -1080 -12080
rect -1000 -12160 -980 -12080
rect -1100 -12180 -980 -12160
rect -600 -11980 -580 -11880
rect -480 -11980 -460 -11880
rect -600 -12000 -460 -11980
rect -600 -12100 -580 -12000
rect -480 -12100 -460 -12000
rect 4440 -11800 4902 -11700
rect 4440 -12100 4560 -11800
rect 4946 -11840 5034 -11540
rect 5640 -11300 5760 -11246
rect 5640 -11340 5860 -11300
rect 5640 -11400 5660 -11340
rect 5720 -11400 5780 -11340
rect 5840 -11400 5860 -11340
rect 5640 -11440 5860 -11400
rect 6100 -11340 6780 -11300
rect 6100 -11400 6160 -11340
rect 6220 -11400 6280 -11340
rect 6340 -11400 6400 -11340
rect 6480 -11400 6540 -11340
rect 6600 -11400 6660 -11340
rect 6720 -11400 6780 -11340
rect 4894 -11902 5034 -11840
rect 5300 -11720 5440 -11700
rect 5300 -11820 5320 -11720
rect 5420 -11820 5440 -11720
rect 5300 -11840 5440 -11820
rect 5300 -11940 5320 -11840
rect 5420 -11940 5440 -11840
rect 5300 -11980 5440 -11940
rect 5300 -12100 5320 -11980
rect 5420 -12100 5440 -11980
rect -600 -12120 -460 -12100
rect -2600 -12580 -2580 -12500
rect -2500 -12580 -2300 -12500
rect -2220 -12580 -2200 -12500
rect -2600 -12600 -2200 -12580
rect -600 -12220 -580 -12120
rect -480 -12220 -460 -12120
rect -600 -12260 -460 -12220
rect -600 -12360 -580 -12260
rect -480 -12360 -460 -12260
rect -600 -12420 -460 -12360
rect -80 -12280 5220 -12100
rect -80 -12284 2320 -12280
rect 2880 -12284 5220 -12280
rect -80 -12420 100 -12284
rect -600 -12600 100 -12420
rect 5040 -12420 5220 -12284
rect 5300 -12140 5440 -12100
rect 5300 -12240 5320 -12140
rect 5420 -12240 5440 -12140
rect 5300 -12260 5440 -12240
rect 5300 -12360 5320 -12260
rect 5420 -12360 5440 -12260
rect 5300 -12380 5440 -12360
rect 5640 -12380 5760 -11440
rect 6100 -11660 6780 -11400
rect 6200 -11700 6760 -11660
rect 6140 -11940 6260 -11920
rect 6140 -12020 6160 -11940
rect 6240 -12020 6260 -11940
rect 6140 -12080 6260 -12020
rect 6140 -12160 6160 -12080
rect 6240 -12160 6260 -12080
rect 6140 -12180 6260 -12160
rect 6720 -11940 6840 -11920
rect 6720 -12020 6740 -11940
rect 6820 -12020 6840 -11940
rect 6720 -12080 6840 -12020
rect 6720 -12160 6740 -12080
rect 6820 -12160 6840 -12080
rect 6720 -12180 6840 -12160
rect 7400 -12020 7800 -12000
rect 7400 -12100 7420 -12020
rect 7500 -12100 7700 -12020
rect 7780 -12100 7800 -12020
rect -600 -12602 -460 -12600
rect 1240 -12880 2140 -12460
rect 2460 -12880 3360 -12460
rect 3660 -12800 3940 -12460
rect 5040 -12600 5640 -12420
rect 7400 -12500 7800 -12100
rect 7400 -12580 7420 -12500
rect 7500 -12580 7700 -12500
rect 7780 -12580 7800 -12500
rect 7400 -12600 7800 -12580
rect 3660 -12860 3700 -12800
rect 3760 -12860 3940 -12800
rect 3660 -12880 3940 -12860
rect 800 -13620 1540 -13500
rect 800 -13680 900 -13620
rect 960 -13680 1540 -13620
rect 800 -13740 1540 -13680
rect 800 -13800 900 -13740
rect 960 -13800 1540 -13740
rect 800 -13920 1540 -13800
rect 800 -14020 1180 -13920
rect 1860 -13940 2760 -13520
rect 3060 -13940 3960 -13520
rect 4020 -14020 4400 -13500
rect 800 -14140 4400 -14020
rect 800 -14200 900 -14140
rect 960 -14200 4400 -14140
rect 800 -14240 4400 -14200
rect 800 -14300 900 -14240
rect 960 -14300 4240 -14240
rect 4300 -14300 4400 -14240
rect 800 -14400 4400 -14300
rect 820 -14680 1080 -14660
rect 820 -14740 840 -14680
rect 900 -14740 1000 -14680
rect 1060 -14740 1080 -14680
rect 820 -14780 1080 -14740
rect 820 -14840 840 -14780
rect 900 -14840 1000 -14780
rect 1060 -14840 1080 -14780
rect 820 -14860 1080 -14840
rect 4120 -14680 4380 -14660
rect 4120 -14740 4140 -14680
rect 4200 -14740 4300 -14680
rect 4360 -14740 4380 -14680
rect 4120 -14780 4380 -14740
rect 4120 -14840 4140 -14780
rect 4200 -14840 4300 -14780
rect 4360 -14840 4380 -14780
rect 4120 -14860 4380 -14840
<< via1 >>
rect 2540 -8560 2620 -8480
rect 2540 -8660 2620 -8580
rect 2540 -8780 2620 -8700
rect 2540 -8880 2620 -8800
rect 2540 -8980 2620 -8900
rect 2540 -9080 2620 -9000
rect 2540 -9180 2620 -9100
rect -1780 -9500 -1700 -9420
rect -1780 -9640 -1700 -9560
rect -1160 -9500 -1080 -9420
rect -1160 -9640 -1080 -9560
rect -540 -9500 -460 -9420
rect -540 -9640 -460 -9560
rect 60 -9500 140 -9420
rect 60 -9640 140 -9560
rect 660 -9500 740 -9420
rect 660 -9640 740 -9560
rect 1780 -9540 1840 -9480
rect 2540 -9280 2620 -9200
rect 2540 -9380 2620 -9300
rect 2360 -9540 2420 -9480
rect 2740 -9540 2800 -9480
rect 3340 -9540 3400 -9480
rect 3960 -9540 4020 -9480
rect 4460 -9500 4540 -9420
rect 4460 -9640 4540 -9560
rect 5040 -9500 5120 -9420
rect 5040 -9640 5120 -9560
rect 5660 -9500 5740 -9420
rect 5660 -9640 5740 -9560
rect 6280 -9500 6360 -9420
rect 6280 -9640 6360 -9560
rect 6880 -9500 6960 -9420
rect 6880 -9640 6960 -9560
rect -3380 -10020 -3300 -9940
rect -3100 -10020 -3020 -9940
rect 3300 -10000 3360 -9940
rect 8220 -10020 8300 -9940
rect 8500 -10020 8580 -9940
rect 3300 -10080 3360 -10020
rect -3380 -10180 -3300 -10100
rect -3100 -10180 -3020 -10100
rect 3300 -10220 3360 -10160
rect 8220 -10180 8300 -10100
rect 8500 -10180 8580 -10100
rect 3300 -10300 3360 -10240
rect -580 -10560 -480 -10460
rect -3540 -10680 -3460 -10600
rect -3540 -10820 -3460 -10740
rect -2960 -10680 -2880 -10600
rect -2960 -10820 -2880 -10740
rect -2340 -10680 -2260 -10600
rect -2340 -10820 -2260 -10740
rect -1720 -10680 -1640 -10600
rect -1720 -10820 -1640 -10740
rect -1140 -10680 -1060 -10600
rect -1140 -10820 -1060 -10740
rect -580 -10760 -480 -10660
rect -580 -10960 -480 -10860
rect 40 -10760 140 -10660
rect 640 -10760 740 -10660
rect 1780 -10480 1840 -10420
rect 2140 -10440 2200 -10380
rect 2240 -10440 2300 -10380
rect 2380 -10440 2440 -10380
rect 2520 -10440 2580 -10380
rect 2620 -10440 2680 -10380
rect 2520 -10540 2580 -10480
rect 2620 -10540 2680 -10480
rect 2760 -10440 2820 -10380
rect 2900 -10440 2960 -10380
rect 3000 -10440 3060 -10380
rect 1780 -10840 1840 -10780
rect 2340 -10840 2400 -10780
rect 2580 -10680 2640 -10620
rect 2820 -10840 2880 -10780
rect 1800 -11000 1860 -10940
rect 3280 -11000 3340 -10940
rect 6240 -10680 6320 -10600
rect 6240 -10820 6320 -10740
rect 6840 -10680 6920 -10600
rect 6840 -10820 6920 -10740
rect 7460 -10680 7540 -10600
rect 7460 -10820 7540 -10740
rect 8080 -10680 8160 -10600
rect 8080 -10820 8160 -10740
rect 8640 -10680 8720 -10600
rect 8640 -10820 8720 -10740
rect 40 -11400 100 -11340
rect 200 -11400 260 -11340
rect 2260 -11660 2320 -11600
rect -580 -11840 -480 -11740
rect 2260 -11760 2320 -11700
rect 2880 -11660 2940 -11600
rect 2880 -11760 2940 -11700
rect -2580 -12100 -2500 -12020
rect -2300 -12100 -2220 -12020
rect -1680 -12020 -1600 -11940
rect -1680 -12160 -1600 -12080
rect -1080 -12020 -1000 -11940
rect -1080 -12160 -1000 -12080
rect -580 -11980 -480 -11880
rect -580 -12100 -480 -12000
rect 5660 -11400 5720 -11340
rect 5780 -11400 5840 -11340
rect 6160 -11400 6220 -11340
rect 6280 -11400 6340 -11340
rect 6400 -11400 6480 -11340
rect 6540 -11400 6600 -11340
rect 6660 -11400 6720 -11340
rect 5320 -11820 5420 -11720
rect 5320 -11940 5420 -11840
rect 5320 -12100 5420 -11980
rect -2580 -12580 -2500 -12500
rect -2300 -12580 -2220 -12500
rect -580 -12220 -480 -12120
rect -580 -12360 -480 -12260
rect 5320 -12240 5420 -12140
rect 5320 -12360 5420 -12260
rect 6160 -12020 6240 -11940
rect 6160 -12160 6240 -12080
rect 6740 -12020 6820 -11940
rect 6740 -12160 6820 -12080
rect 7420 -12100 7500 -12020
rect 7700 -12100 7780 -12020
rect 7420 -12580 7500 -12500
rect 7700 -12580 7780 -12500
rect 3700 -12860 3760 -12800
rect 840 -14740 900 -14680
rect 1000 -14740 1060 -14680
rect 840 -14840 900 -14780
rect 1000 -14840 1060 -14780
rect 4140 -14740 4200 -14680
rect 4300 -14740 4360 -14680
rect 4140 -14840 4200 -14780
rect 4300 -14840 4360 -14780
<< metal2 >>
rect 2500 -8480 2660 -8460
rect 2500 -8560 2540 -8480
rect 2620 -8560 2660 -8480
rect 2500 -8580 2660 -8560
rect 2500 -8660 2540 -8580
rect 2620 -8660 2660 -8580
rect 2500 -8700 2660 -8660
rect 2500 -8780 2540 -8700
rect 2620 -8780 2660 -8700
rect 2500 -8800 2660 -8780
rect 2500 -8880 2540 -8800
rect 2620 -8880 2660 -8800
rect 2500 -8900 2660 -8880
rect 2500 -8980 2540 -8900
rect 2620 -8980 2660 -8900
rect 2500 -9000 2660 -8980
rect 2500 -9080 2540 -9000
rect 2620 -9080 2660 -9000
rect 2500 -9100 2660 -9080
rect 2500 -9140 2540 -9100
rect 360 -9180 2540 -9140
rect 2620 -9140 2660 -9100
rect 2620 -9180 4840 -9140
rect 360 -9200 4840 -9180
rect 360 -9280 2540 -9200
rect 2620 -9280 4840 -9200
rect 360 -9300 4840 -9280
rect 360 -9380 2540 -9300
rect 2620 -9380 4840 -9300
rect 360 -9400 4840 -9380
rect -2140 -9420 760 -9400
rect -2140 -9500 -1780 -9420
rect -1700 -9500 -1160 -9420
rect -1080 -9500 -540 -9420
rect -460 -9500 60 -9420
rect 140 -9500 660 -9420
rect 740 -9500 760 -9420
rect 4440 -9420 7340 -9400
rect -2140 -9560 760 -9500
rect -3400 -9940 -3000 -9600
rect -3400 -10020 -3380 -9940
rect -3300 -10020 -3100 -9940
rect -3020 -10020 -3000 -9940
rect -3400 -10100 -3000 -10020
rect -3400 -10180 -3380 -10100
rect -3300 -10180 -3100 -10100
rect -3020 -10180 -3000 -10100
rect -3400 -10200 -3000 -10180
rect -2140 -9640 -1780 -9560
rect -1700 -9640 -1160 -9560
rect -1080 -9640 -540 -9560
rect -460 -9640 60 -9560
rect 140 -9640 660 -9560
rect 740 -9640 760 -9560
rect 1120 -9480 2460 -9440
rect 1120 -9540 1780 -9480
rect 1840 -9540 2360 -9480
rect 2420 -9540 2460 -9480
rect 1120 -9580 2460 -9540
rect 2720 -9480 4040 -9440
rect 2720 -9540 2740 -9480
rect 2800 -9540 3340 -9480
rect 3400 -9540 3960 -9480
rect 4020 -9540 4040 -9480
rect 2720 -9580 4040 -9540
rect 4440 -9500 4460 -9420
rect 4540 -9500 5040 -9420
rect 5120 -9500 5660 -9420
rect 5740 -9500 6280 -9420
rect 6360 -9500 6880 -9420
rect 6960 -9500 7340 -9420
rect 4440 -9560 7340 -9500
rect -2140 -9660 760 -9640
rect -2140 -10580 -1840 -9660
rect 1760 -10420 1860 -9580
rect 3280 -9940 3380 -9580
rect 4440 -9640 4460 -9560
rect 4540 -9640 5040 -9560
rect 5120 -9640 5660 -9560
rect 5740 -9640 6280 -9560
rect 6360 -9640 6880 -9560
rect 6960 -9640 7340 -9560
rect 4440 -9660 7340 -9640
rect 3280 -10000 3300 -9940
rect 3360 -10000 3380 -9940
rect 3280 -10020 3380 -10000
rect 3280 -10080 3300 -10020
rect 3360 -10080 3380 -10020
rect 3280 -10160 3380 -10080
rect 2460 -10200 2740 -10180
rect 2460 -10260 2480 -10200
rect 2540 -10260 2660 -10200
rect 2720 -10260 2740 -10200
rect 2460 -10280 2740 -10260
rect 3280 -10220 3300 -10160
rect 3360 -10220 3380 -10160
rect 3280 -10240 3380 -10220
rect 3280 -10300 3300 -10240
rect 3360 -10300 3380 -10240
rect -600 -10460 -460 -10440
rect -600 -10560 -580 -10460
rect -480 -10560 -460 -10460
rect 1760 -10480 1780 -10420
rect 1840 -10480 1860 -10420
rect 2120 -10380 2460 -10360
rect 2120 -10440 2140 -10380
rect 2200 -10440 2240 -10380
rect 2300 -10440 2380 -10380
rect 2440 -10440 2460 -10380
rect 2120 -10460 2460 -10440
rect 2500 -10380 2700 -10360
rect 2500 -10440 2520 -10380
rect 2580 -10440 2620 -10380
rect 2680 -10440 2700 -10380
rect 1760 -10500 1860 -10480
rect 2500 -10480 2700 -10440
rect 2740 -10380 3080 -10360
rect 2740 -10440 2760 -10380
rect 2820 -10440 2900 -10380
rect 2960 -10440 3000 -10380
rect 3060 -10440 3080 -10380
rect 2740 -10460 3080 -10440
rect 2500 -10540 2520 -10480
rect 2580 -10540 2620 -10480
rect 2680 -10540 2700 -10480
rect 2500 -10560 2700 -10540
rect -3560 -10600 -1040 -10580
rect -3560 -10680 -3540 -10600
rect -3460 -10680 -2960 -10600
rect -2880 -10680 -2340 -10600
rect -2260 -10680 -1720 -10600
rect -1640 -10680 -1140 -10600
rect -1060 -10680 -1040 -10600
rect -3560 -10740 -1040 -10680
rect -3560 -10820 -3540 -10740
rect -3460 -10820 -2960 -10740
rect -2880 -10820 -2340 -10740
rect -2260 -10820 -1720 -10740
rect -1640 -10820 -1140 -10740
rect -1060 -10820 -1040 -10740
rect -3560 -10840 -1040 -10820
rect -600 -10640 -460 -10560
rect 3280 -10600 3380 -10300
rect 7040 -10580 7340 -9660
rect 8200 -9940 8600 -9600
rect 8200 -10020 8220 -9940
rect 8300 -10020 8500 -9940
rect 8580 -10020 8600 -9940
rect 8200 -10100 8600 -10020
rect 8200 -10180 8220 -10100
rect 8300 -10180 8500 -10100
rect 8580 -10180 8600 -10100
rect 8200 -10200 8600 -10180
rect 1760 -10620 3380 -10600
rect -600 -10660 760 -10640
rect -600 -10760 -580 -10660
rect -480 -10760 40 -10660
rect 140 -10760 640 -10660
rect 740 -10760 760 -10660
rect 1760 -10680 2580 -10620
rect 2640 -10680 3380 -10620
rect 1760 -10700 3380 -10680
rect 6220 -10600 8740 -10580
rect 6220 -10680 6240 -10600
rect 6320 -10680 6840 -10600
rect 6920 -10680 7460 -10600
rect 7540 -10680 8080 -10600
rect 8160 -10680 8640 -10600
rect 8720 -10680 8740 -10600
rect 6220 -10740 8740 -10680
rect -600 -10780 760 -10760
rect 1760 -10780 3380 -10760
rect -2140 -11920 -1840 -10840
rect -600 -10860 -460 -10780
rect 1760 -10840 1780 -10780
rect 1840 -10840 2340 -10780
rect 2400 -10840 2820 -10780
rect 2880 -10840 3380 -10780
rect 6220 -10820 6240 -10740
rect 6320 -10820 6840 -10740
rect 6920 -10820 7460 -10740
rect 7540 -10820 8080 -10740
rect 8160 -10820 8640 -10740
rect 8720 -10820 8740 -10740
rect 6220 -10840 8740 -10820
rect 1760 -10860 3380 -10840
rect -600 -10960 -580 -10860
rect -480 -10960 -460 -10860
rect -1640 -11340 -960 -11300
rect -1640 -11400 -1580 -11340
rect -1520 -11400 -1460 -11340
rect -1400 -11400 -1340 -11340
rect -1260 -11400 -1200 -11340
rect -1140 -11400 -1080 -11340
rect -1020 -11400 -960 -11340
rect -1640 -11440 -960 -11400
rect -600 -11740 -460 -10960
rect 1760 -10940 1900 -10920
rect 1760 -11000 1800 -10940
rect 1860 -11000 1900 -10940
rect -360 -11340 280 -11300
rect -360 -11400 -340 -11340
rect -280 -11400 -220 -11340
rect -160 -11400 40 -11340
rect 100 -11400 200 -11340
rect 260 -11400 280 -11340
rect -360 -11440 280 -11400
rect -600 -11840 -580 -11740
rect -480 -11840 -460 -11740
rect 1760 -11580 1900 -11000
rect 3240 -10940 3380 -10920
rect 3240 -11000 3280 -10940
rect 3340 -11000 3380 -10940
rect 3240 -11580 3380 -11000
rect 5640 -11340 6780 -11300
rect 5640 -11400 5660 -11340
rect 5720 -11400 5780 -11340
rect 5840 -11400 6160 -11340
rect 6220 -11400 6280 -11340
rect 6340 -11400 6400 -11340
rect 6480 -11400 6540 -11340
rect 6600 -11400 6660 -11340
rect 6720 -11400 6780 -11340
rect 5640 -11440 6780 -11400
rect 1760 -11600 3380 -11580
rect 1760 -11660 2260 -11600
rect 2320 -11660 2880 -11600
rect 2940 -11660 3380 -11600
rect 1760 -11700 3380 -11660
rect 1760 -11760 2260 -11700
rect 2320 -11760 2880 -11700
rect 2940 -11760 3380 -11700
rect 1760 -11780 3380 -11760
rect 5300 -11720 5440 -11700
rect -600 -11880 -460 -11840
rect -2540 -11940 -980 -11920
rect -2540 -12000 -1680 -11940
rect -2600 -12020 -1680 -12000
rect -1600 -12020 -1080 -11940
rect -1000 -12020 -980 -11940
rect -2600 -12100 -2580 -12020
rect -2500 -12100 -2300 -12020
rect -2220 -12080 -980 -12020
rect -2220 -12100 -1680 -12080
rect -2600 -12160 -1680 -12100
rect -1600 -12160 -1080 -12080
rect -1000 -12160 -980 -12080
rect -2600 -12180 -980 -12160
rect -600 -11980 -580 -11880
rect -480 -11980 -460 -11880
rect -600 -12000 -460 -11980
rect -600 -12100 -580 -12000
rect -480 -12100 -460 -12000
rect -600 -12120 -460 -12100
rect -2600 -12500 -2200 -12180
rect -600 -12220 -580 -12120
rect -480 -12220 -460 -12120
rect -600 -12260 -460 -12220
rect -600 -12360 -580 -12260
rect -480 -12360 -460 -12260
rect -600 -12380 -460 -12360
rect 5300 -11820 5320 -11720
rect 5420 -11820 5440 -11720
rect 5300 -11840 5440 -11820
rect 5300 -11940 5320 -11840
rect 5420 -11940 5440 -11840
rect 7040 -11920 7340 -10840
rect 5300 -11980 5440 -11940
rect 5300 -12100 5320 -11980
rect 5420 -12100 5440 -11980
rect 5300 -12140 5440 -12100
rect 5300 -12240 5320 -12140
rect 5420 -12240 5440 -12140
rect 6140 -11940 7700 -11920
rect 6140 -12020 6160 -11940
rect 6240 -12020 6740 -11940
rect 6820 -12000 7700 -11940
rect 6820 -12020 7800 -12000
rect 6140 -12080 7420 -12020
rect 6140 -12160 6160 -12080
rect 6240 -12160 6740 -12080
rect 6820 -12100 7420 -12080
rect 7500 -12100 7700 -12020
rect 7780 -12100 7800 -12020
rect 6820 -12160 7800 -12100
rect 6140 -12180 7800 -12160
rect 5300 -12260 5440 -12240
rect 5300 -12360 5320 -12260
rect 5420 -12360 5440 -12260
rect 5300 -12440 5440 -12360
rect -2600 -12580 -2580 -12500
rect -2500 -12580 -2300 -12500
rect -2220 -12580 -2200 -12500
rect -2600 -12600 -2200 -12580
rect 3660 -12800 5480 -12440
rect 7400 -12500 7800 -12180
rect 7400 -12580 7420 -12500
rect 7500 -12580 7700 -12500
rect 7780 -12580 7800 -12500
rect 7400 -12600 7800 -12580
rect 3660 -12860 3700 -12800
rect 3760 -12860 5480 -12800
rect 3660 -12880 5480 -12860
rect 5300 -12900 5440 -12880
rect 820 -14680 1080 -14660
rect 820 -14740 840 -14680
rect 900 -14740 1000 -14680
rect 1060 -14740 1080 -14680
rect 820 -14780 1080 -14740
rect 820 -14840 840 -14780
rect 900 -14840 1000 -14780
rect 1060 -14840 1080 -14780
rect 820 -14860 1080 -14840
rect 4120 -14680 4380 -14660
rect 4120 -14740 4140 -14680
rect 4200 -14740 4300 -14680
rect 4360 -14740 4380 -14680
rect 4120 -14780 4380 -14740
rect 4120 -14840 4140 -14780
rect 4200 -14840 4300 -14780
rect 4360 -14840 4380 -14780
rect 4120 -14860 4380 -14840
<< via2 >>
rect -3380 -10020 -3300 -9940
rect -3100 -10020 -3020 -9940
rect -3380 -10180 -3300 -10100
rect -3100 -10180 -3020 -10100
rect 2480 -10260 2540 -10200
rect 2660 -10260 2720 -10200
rect 2140 -10440 2200 -10380
rect 2240 -10440 2300 -10380
rect 2520 -10440 2580 -10380
rect 2620 -10440 2680 -10380
rect 2900 -10440 2960 -10380
rect 3000 -10440 3060 -10380
rect 2520 -10540 2580 -10480
rect 2620 -10540 2680 -10480
rect 8220 -10020 8300 -9940
rect 8500 -10020 8580 -9940
rect 8220 -10180 8300 -10100
rect 8500 -10180 8580 -10100
rect -1580 -11400 -1520 -11340
rect -1460 -11400 -1400 -11340
rect -1340 -11400 -1260 -11340
rect -1200 -11400 -1140 -11340
rect -1080 -11400 -1020 -11340
rect -340 -11400 -280 -11340
rect -220 -11400 -160 -11340
rect -2580 -12100 -2500 -12020
rect -2300 -12100 -2220 -12020
rect 7420 -12100 7500 -12020
rect 7700 -12100 7780 -12020
rect -2580 -12580 -2500 -12500
rect -2300 -12580 -2220 -12500
rect 7420 -12580 7500 -12500
rect 7700 -12580 7780 -12500
rect 840 -14740 900 -14680
rect 1000 -14740 1060 -14680
rect 840 -14840 900 -14780
rect 1000 -14840 1060 -14780
rect 4140 -14740 4200 -14680
rect 4300 -14740 4360 -14680
rect 4140 -14840 4200 -14780
rect 4300 -14840 4360 -14780
<< metal3 >>
rect -3400 -9940 -3000 -9600
rect -3400 -10020 -3380 -9940
rect -3300 -10020 -3100 -9940
rect -3020 -10020 -3000 -9940
rect -3400 -10100 -3000 -10020
rect -3400 -10180 -3380 -10100
rect -3300 -10180 -3100 -10100
rect -3020 -10180 -3000 -10100
rect 8200 -9940 8600 -9600
rect 8200 -10020 8220 -9940
rect 8300 -10020 8500 -9940
rect 8580 -10020 8600 -9940
rect 8200 -10100 8600 -10020
rect 8200 -10180 8220 -10100
rect 8300 -10180 8500 -10100
rect 8580 -10180 8600 -10100
rect -3400 -10200 -3000 -10180
rect 820 -10200 4380 -10180
rect 8200 -10200 8600 -10180
rect 820 -10260 2480 -10200
rect 2540 -10260 2660 -10200
rect 2720 -10260 4380 -10200
rect 820 -10280 4380 -10260
rect 2120 -10360 2420 -10340
rect 820 -10440 2140 -10360
rect 2220 -10380 2320 -10360
rect 2220 -10440 2240 -10380
rect 2300 -10440 2320 -10380
rect 2400 -10440 2420 -10360
rect 820 -10460 2420 -10440
rect 2500 -10380 2700 -10280
rect 2500 -10440 2520 -10380
rect 2580 -10440 2620 -10380
rect 2680 -10440 2700 -10380
rect -1640 -11340 -140 -11300
rect -1640 -11400 -1580 -11340
rect -1520 -11400 -1460 -11340
rect -1400 -11400 -1340 -11340
rect -1260 -11400 -1200 -11340
rect -1140 -11400 -1080 -11340
rect -1020 -11400 -340 -11340
rect -280 -11400 -220 -11340
rect -160 -11400 -140 -11340
rect -1640 -11440 -140 -11400
rect -2600 -12020 -2200 -12000
rect -2600 -12100 -2580 -12020
rect -2500 -12100 -2300 -12020
rect -2220 -12100 -2200 -12020
rect -2600 -12500 -2200 -12100
rect -2600 -12580 -2580 -12500
rect -2500 -12580 -2300 -12500
rect -2220 -12580 -2200 -12500
rect -2600 -12600 -2200 -12580
rect 820 -14680 1080 -10460
rect 2500 -10480 2700 -10440
rect 2780 -10360 3080 -10340
rect 2780 -10440 2800 -10360
rect 2880 -10380 2980 -10360
rect 2880 -10440 2900 -10380
rect 2960 -10440 2980 -10380
rect 3060 -10440 3740 -10360
rect 2780 -10460 3740 -10440
rect 2500 -10540 2520 -10480
rect 2580 -10540 2620 -10480
rect 2680 -10540 2700 -10480
rect 2500 -10560 2700 -10540
rect 820 -14740 840 -14680
rect 900 -14740 1000 -14680
rect 1060 -14740 1080 -14680
rect 820 -14780 1080 -14740
rect 820 -14840 840 -14780
rect 900 -14840 1000 -14780
rect 1060 -14840 1080 -14780
rect 820 -14860 1080 -14840
rect 4120 -14680 4380 -10280
rect 7400 -12020 7800 -12000
rect 7400 -12100 7420 -12020
rect 7500 -12100 7700 -12020
rect 7780 -12100 7800 -12020
rect 7400 -12500 7800 -12100
rect 7400 -12580 7420 -12500
rect 7500 -12580 7700 -12500
rect 7780 -12580 7800 -12500
rect 7400 -12600 7800 -12580
rect 4120 -14740 4140 -14680
rect 4200 -14740 4300 -14680
rect 4360 -14740 4380 -14680
rect 4120 -14780 4380 -14740
rect 4120 -14840 4140 -14780
rect 4200 -14840 4300 -14780
rect 4360 -14840 4380 -14780
rect 4120 -14860 4380 -14840
<< via3 >>
rect -3380 -10020 -3300 -9940
rect -3100 -10020 -3020 -9940
rect -3380 -10180 -3300 -10100
rect -3100 -10180 -3020 -10100
rect 8220 -10020 8300 -9940
rect 8500 -10020 8580 -9940
rect 8220 -10180 8300 -10100
rect 8500 -10180 8580 -10100
rect 2140 -10380 2220 -10360
rect 2140 -10440 2200 -10380
rect 2200 -10440 2220 -10380
rect 2320 -10440 2400 -10360
rect -2580 -12100 -2500 -12020
rect -2300 -12100 -2220 -12020
rect -2580 -12580 -2500 -12500
rect -2300 -12580 -2220 -12500
rect 2800 -10440 2880 -10360
rect 2980 -10380 3060 -10360
rect 2980 -10440 3000 -10380
rect 3000 -10440 3060 -10380
rect 7420 -12100 7500 -12020
rect 7700 -12100 7780 -12020
rect 7420 -12580 7500 -12500
rect 7700 -12580 7780 -12500
<< metal4 >>
rect -6200 -15200 -5800 -8200
rect -4400 -8600 9600 -8200
rect -4400 -15000 -4000 -8600
rect -3400 -9940 -3000 -8600
rect -3400 -10020 -3380 -9940
rect -3300 -10020 -3100 -9940
rect -3020 -10020 -3000 -9940
rect -3400 -10100 -3000 -10020
rect -3400 -10180 -3380 -10100
rect -3300 -10180 -3100 -10100
rect -3020 -10180 -3000 -10100
rect -3400 -10200 -3000 -10180
rect 8200 -9940 8600 -8600
rect 8200 -10020 8220 -9940
rect 8300 -10020 8500 -9940
rect 8580 -10020 8600 -9940
rect 8200 -10100 8600 -10020
rect 8200 -10180 8220 -10100
rect 8300 -10180 8500 -10100
rect 8580 -10180 8600 -10100
rect 8200 -10200 8600 -10180
rect 2120 -10360 2420 -10340
rect 2780 -10360 3080 -10340
rect 2120 -10440 2140 -10360
rect 2220 -10440 2320 -10360
rect 2400 -10440 2800 -10360
rect 2880 -10440 2980 -10360
rect 3060 -10440 3080 -10360
rect 2120 -10460 3080 -10440
rect -2600 -12020 -2200 -12000
rect -2600 -12100 -2580 -12020
rect -2500 -12100 -2300 -12020
rect -2220 -12100 -2200 -12020
rect -2600 -12500 -2200 -12100
rect -2600 -12580 -2580 -12500
rect -2500 -12580 -2300 -12500
rect -2220 -12580 -2200 -12500
rect -2600 -15200 -2200 -12580
rect 7400 -12020 7800 -12000
rect 7400 -12100 7420 -12020
rect 7500 -12100 7700 -12020
rect 7780 -12100 7800 -12020
rect 7400 -12500 7800 -12100
rect 7400 -12580 7420 -12500
rect 7500 -12580 7700 -12500
rect 7780 -12580 7800 -12500
rect 7400 -15200 7800 -12580
rect 9200 -15000 9600 -8600
rect 11000 -15200 11400 -8200
rect -6200 -15600 11400 -15200
use sky130_fd_pr__cap_mim_m3_1_HGL9NV  sky130_fd_pr__cap_mim_m3_1_HGL9NV_0
timestamp 1771116256
transform 1 0 -5914 0 1 -11680
box -1686 -3320 1686 3320
use sky130_fd_pr__nfet_01v8_P5W7CC  sky130_fd_pr__nfet_01v8_P5W7CC_0
timestamp 1771126488
transform 1 0 -1325 0 1 -12021
box -475 -479 475 479
use sky130_fd_pr__nfet_01v8_RJXUD9  sky130_fd_pr__nfet_01v8_RJXUD9_0
timestamp 1771119226
transform 1 0 -379 0 1 -12081
box -321 -519 321 519
use sky130_fd_pr__pfet_01v8_55LJLG  sky130_fd_pr__pfet_01v8_55LJLG_0
timestamp 1771116256
transform 1 0 7499 0 1 -10672
box -1399 -528 1399 528
use sky130_fd_pr__pfet_01v8_55LJLG  sky130_fd_pr__pfet_01v8_55LJLG_1
timestamp 1771116256
transform 1 0 -2301 0 1 -10672
box -1399 -528 1399 528
use sky130_fd_pr__pfet_01v8_EAP5WJ  sky130_fd_pr__pfet_01v8_EAP5WJ_0
timestamp 1771119226
transform 1 0 1783 0 1 -9546
box -783 -454 783 454
use sky130_fd_pr__pfet_01v8_JEJJ38  sky130_fd_pr__pfet_01v8_JEJJ38_0
timestamp 1771116256
transform 1 0 5699 0 1 -9572
box -1399 -528 1399 528
use sky130_fd_pr__pfet_01v8_JEJJ38  sky130_fd_pr__pfet_01v8_JEJJ38_1
timestamp 1771116256
transform 1 0 -501 0 1 -9572
box -1399 -528 1399 528
use sky130_fd_pr__cap_mim_m3_1_HGL9NV  XC2
timestamp 1771116256
transform -1 0 11086 0 -1 -11680
box -1686 -3320 1686 3320
use sky130_fd_pr__nfet_01v8_CSRU6X  XM1
timestamp 1771117290
transform 1 0 2603 0 1 -10696
box -403 -304 403 304
use sky130_fd_pr__pfet_01v8_EAP5WJ  XM3
timestamp 1771119226
transform 1 0 3383 0 1 -9546
box -783 -454 783 454
use sky130_fd_pr__nfet_01v8_6UV5Z4  XM5
timestamp 1771126488
transform 1 0 2595 0 1 -11681
box -475 -519 475 519
use sky130_fd_pr__nfet_01v8_P5W7CC  XM7
timestamp 1771126488
transform 1 0 6475 0 1 -12021
box -475 -479 475 479
use sky130_fd_pr__pfet_01v8_EAP5WJ  XM8
timestamp 1771119226
transform 1 0 5083 0 1 -10746
box -783 -454 783 454
use sky130_fd_pr__nfet_01v8_RJXUD9  XM10
timestamp 1771119226
transform 1 0 5521 0 1 -12081
box -321 -519 321 519
use sky130_fd_pr__pfet_01v8_EAP5WJ  XM11
timestamp 1771119226
transform 1 0 83 0 1 -10746
box -783 -454 783 454
use sky130_fd_pr__nfet_01v8_TYFUPF  XM12
timestamp 1771143426
transform 1 0 4927 0 1 -11723
box -211 -295 211 295
use sky130_fd_pr__res_high_po_1p41_B3F3CB  XR2
timestamp 1771116256
transform 1 0 1407 0 1 -13194
box -307 -906 307 906
use sky130_fd_pr__res_high_po_1p41_B3F3CB  XR3
timestamp 1771116256
transform 1 0 2007 0 1 -13194
box -307 -906 307 906
use sky130_fd_pr__res_high_po_1p41_B3F3CB  XR4
timestamp 1771116256
transform 1 0 2607 0 1 -13194
box -307 -906 307 906
use sky130_fd_pr__res_high_po_1p41_B3F3CB  XR5
timestamp 1771116256
transform 1 0 3207 0 1 -13194
box -307 -906 307 906
use sky130_fd_pr__res_high_po_1p41_B3F3CB  XR6
timestamp 1771116256
transform 1 0 3807 0 1 -13194
box -307 -906 307 906
<< labels >>
flabel metal1 880 -13800 1080 -13600 0 FreeSans 256 0 0 0 VSS
port 4 nsew
flabel metal1 2480 -8660 2680 -8460 0 FreeSans 256 0 0 0 OUT
port 1 nsew
flabel locali -3380 -9440 -3180 -9240 0 FreeSans 1600 0 0 0 VDD
port 6 nsew
flabel metal1 880 -14860 1080 -14660 0 FreeSans 256 0 0 0 VP
port 2 nsew
flabel metal1 4120 -14860 4320 -14660 0 FreeSans 256 0 0 0 VN
port 3 nsew
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1770979109
<< xpolycontact >>
rect -141 125 141 557
rect -141 -557 141 -125
<< xpolyres >>
rect -141 -125 141 125
<< viali >>
rect -125 142 125 539
rect -125 -539 125 -142
<< metal1 >>
rect -131 539 131 551
rect -131 142 -125 539
rect 125 142 131 539
rect -131 130 131 142
rect -131 -142 131 -130
rect -131 -539 -125 -142
rect 125 -539 131 -142
rect -131 -551 131 -539
<< properties >>
string gencell sky130_fd_pr__res_xhigh_po_1p41
string library sky130
string parameters w 1.410 l 1.41 m 1 nx 1 wmin 1.410 lmin 0.50 class resistor rho 2000 val 2.266k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 1.410 guard 0 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1771420802
<< error_p >>
rect -530 3424 530 3436
rect -530 -3424 -518 3424
rect -494 3388 494 3400
rect -494 3284 -482 3388
rect -301 3328 -179 3331
rect -141 3328 -19 3331
rect 19 3328 141 3331
rect 179 3328 301 3331
rect -481 3284 -465 3300
rect -451 3284 -435 3300
rect -263 3293 -247 3309
rect -233 3293 -217 3309
rect -103 3293 -87 3309
rect -73 3293 -57 3309
rect 57 3293 73 3309
rect 87 3293 103 3309
rect 217 3293 233 3309
rect 247 3293 263 3309
rect -497 3268 -481 3284
rect -435 3268 -419 3284
rect -279 3277 -201 3293
rect -119 3277 -41 3293
rect 41 3277 119 3293
rect 201 3277 279 3293
rect 435 3284 451 3300
rect 465 3284 481 3300
rect 482 3284 494 3388
rect -494 -3268 -482 3268
rect -274 3263 -206 3277
rect -114 3263 -46 3277
rect 46 3263 114 3277
rect 206 3263 274 3277
rect 419 3268 435 3284
rect 481 3268 497 3284
rect -279 3247 -201 3263
rect -119 3247 -41 3263
rect 41 3247 119 3263
rect 201 3247 279 3263
rect -263 3231 -247 3247
rect -233 3231 -217 3247
rect -103 3231 -87 3247
rect -73 3231 -57 3247
rect 57 3231 73 3247
rect 87 3231 103 3247
rect 217 3231 233 3247
rect 247 3231 263 3247
rect -343 3201 -327 3217
rect -313 3201 -297 3217
rect -183 3201 -167 3217
rect -153 3201 -137 3217
rect -23 3201 -7 3217
rect 7 3201 23 3217
rect 137 3201 153 3217
rect 167 3201 183 3217
rect 297 3201 313 3217
rect 327 3201 343 3217
rect -359 3185 -343 3201
rect -297 3185 -281 3201
rect -199 3185 -183 3201
rect -137 3185 -121 3201
rect -39 3185 -23 3201
rect 23 3185 39 3201
rect 121 3185 137 3201
rect 183 3185 199 3201
rect 281 3185 297 3201
rect 343 3185 359 3201
rect -359 2127 -343 2143
rect -297 2128 -281 2143
rect -199 2128 -183 2143
rect -297 2127 -183 2128
rect -137 2128 -121 2143
rect -39 2128 -23 2143
rect -137 2127 -23 2128
rect 23 2128 39 2143
rect 121 2128 137 2143
rect 23 2127 137 2128
rect 183 2128 199 2143
rect 281 2128 297 2143
rect 183 2127 297 2128
rect 343 2127 359 2143
rect -343 2111 -327 2127
rect -313 2114 -167 2127
rect -313 2111 -297 2114
rect -183 2111 -167 2114
rect -153 2114 -7 2127
rect -153 2111 -137 2114
rect -23 2111 -7 2114
rect 7 2114 153 2127
rect 7 2111 23 2114
rect 137 2111 153 2114
rect 167 2114 313 2127
rect 167 2111 183 2114
rect 297 2111 313 2114
rect 327 2111 343 2127
rect -263 2081 -247 2097
rect -233 2081 -217 2097
rect -103 2081 -87 2097
rect -73 2081 -57 2097
rect 57 2081 73 2097
rect 87 2081 103 2097
rect 217 2081 233 2097
rect 247 2081 263 2097
rect -279 2065 -201 2081
rect -119 2065 -41 2081
rect 41 2065 119 2081
rect 201 2065 279 2081
rect -274 2051 -206 2065
rect -114 2051 -46 2065
rect 46 2051 114 2065
rect 206 2051 274 2065
rect -279 2035 -201 2051
rect -119 2035 -41 2051
rect 41 2035 119 2051
rect 201 2035 279 2051
rect -263 2019 -247 2035
rect -233 2019 -217 2035
rect -103 2019 -87 2035
rect -73 2019 -57 2035
rect 57 2019 73 2035
rect 87 2019 103 2035
rect 217 2019 233 2035
rect 247 2019 263 2035
rect -263 1961 -247 1977
rect -233 1961 -217 1977
rect -103 1961 -87 1977
rect -73 1961 -57 1977
rect 57 1961 73 1977
rect 87 1961 103 1977
rect 217 1961 233 1977
rect 247 1961 263 1977
rect -279 1945 -201 1961
rect -119 1945 -41 1961
rect 41 1945 119 1961
rect 201 1945 279 1961
rect -274 1931 -206 1945
rect -114 1931 -46 1945
rect 46 1931 114 1945
rect 206 1931 274 1945
rect -279 1915 -201 1931
rect -119 1915 -41 1931
rect 41 1915 119 1931
rect 201 1915 279 1931
rect -263 1899 -247 1915
rect -233 1899 -217 1915
rect -103 1899 -87 1915
rect -73 1899 -57 1915
rect 57 1899 73 1915
rect 87 1899 103 1915
rect 217 1899 233 1915
rect 247 1899 263 1915
rect -343 1869 -327 1885
rect -313 1869 -297 1885
rect -183 1869 -167 1885
rect -153 1869 -137 1885
rect -23 1869 -7 1885
rect 7 1869 23 1885
rect 137 1869 153 1885
rect 167 1869 183 1885
rect 297 1869 313 1885
rect 327 1869 343 1885
rect -359 1853 -343 1869
rect -297 1853 -281 1869
rect -199 1853 -183 1869
rect -137 1853 -121 1869
rect -39 1853 -23 1869
rect 23 1853 39 1869
rect 121 1853 137 1869
rect 183 1853 199 1869
rect 281 1853 297 1869
rect 343 1853 359 1869
rect -359 795 -343 811
rect -297 796 -281 811
rect -199 796 -183 811
rect -297 795 -183 796
rect -137 796 -121 811
rect -39 796 -23 811
rect -137 795 -23 796
rect 23 796 39 811
rect 121 796 137 811
rect 23 795 137 796
rect 183 796 199 811
rect 281 796 297 811
rect 183 795 297 796
rect 343 795 359 811
rect -343 779 -327 795
rect -313 782 -167 795
rect -313 779 -297 782
rect -183 779 -167 782
rect -153 782 -7 795
rect -153 779 -137 782
rect -23 779 -7 782
rect 7 782 153 795
rect 7 779 23 782
rect 137 779 153 782
rect 167 782 313 795
rect 167 779 183 782
rect 297 779 313 782
rect 327 779 343 795
rect -263 749 -247 765
rect -233 749 -217 765
rect -103 749 -87 765
rect -73 749 -57 765
rect 57 749 73 765
rect 87 749 103 765
rect 217 749 233 765
rect 247 749 263 765
rect -279 733 -201 749
rect -119 733 -41 749
rect 41 733 119 749
rect 201 733 279 749
rect -274 719 -206 733
rect -114 719 -46 733
rect 46 719 114 733
rect 206 719 274 733
rect -279 703 -201 719
rect -119 703 -41 719
rect 41 703 119 719
rect 201 703 279 719
rect -263 687 -247 703
rect -233 687 -217 703
rect -103 687 -87 703
rect -73 687 -57 703
rect 57 687 73 703
rect 87 687 103 703
rect 217 687 233 703
rect 247 687 263 703
rect -263 629 -247 645
rect -233 629 -217 645
rect -103 629 -87 645
rect -73 629 -57 645
rect 57 629 73 645
rect 87 629 103 645
rect 217 629 233 645
rect 247 629 263 645
rect -279 613 -201 629
rect -119 613 -41 629
rect 41 613 119 629
rect 201 613 279 629
rect -274 599 -206 613
rect -114 599 -46 613
rect 46 599 114 613
rect 206 599 274 613
rect -279 583 -201 599
rect -119 583 -41 599
rect 41 583 119 599
rect 201 583 279 599
rect -263 567 -247 583
rect -233 567 -217 583
rect -103 567 -87 583
rect -73 567 -57 583
rect 57 567 73 583
rect 87 567 103 583
rect 217 567 233 583
rect 247 567 263 583
rect -343 537 -327 553
rect -313 537 -297 553
rect -183 537 -167 553
rect -153 537 -137 553
rect -23 537 -7 553
rect 7 537 23 553
rect 137 537 153 553
rect 167 537 183 553
rect 297 537 313 553
rect 327 537 343 553
rect -359 521 -343 537
rect -297 521 -281 537
rect -199 521 -183 537
rect -137 521 -121 537
rect -39 521 -23 537
rect 23 521 39 537
rect 121 521 137 537
rect 183 521 199 537
rect 281 521 297 537
rect 343 521 359 537
rect -359 -537 -343 -521
rect -297 -536 -281 -521
rect -199 -536 -183 -521
rect -297 -537 -183 -536
rect -137 -536 -121 -521
rect -39 -536 -23 -521
rect -137 -537 -23 -536
rect 23 -536 39 -521
rect 121 -536 137 -521
rect 23 -537 137 -536
rect 183 -536 199 -521
rect 281 -536 297 -521
rect 183 -537 297 -536
rect 343 -537 359 -521
rect -343 -553 -327 -537
rect -313 -550 -167 -537
rect -313 -553 -297 -550
rect -183 -553 -167 -550
rect -153 -550 -7 -537
rect -153 -553 -137 -550
rect -23 -553 -7 -550
rect 7 -550 153 -537
rect 7 -553 23 -550
rect 137 -553 153 -550
rect 167 -550 313 -537
rect 167 -553 183 -550
rect 297 -553 313 -550
rect 327 -553 343 -537
rect -263 -583 -247 -567
rect -233 -583 -217 -567
rect -103 -583 -87 -567
rect -73 -583 -57 -567
rect 57 -583 73 -567
rect 87 -583 103 -567
rect 217 -583 233 -567
rect 247 -583 263 -567
rect -279 -599 -201 -583
rect -119 -599 -41 -583
rect 41 -599 119 -583
rect 201 -599 279 -583
rect -274 -613 -206 -599
rect -114 -613 -46 -599
rect 46 -613 114 -599
rect 206 -613 274 -599
rect -279 -629 -201 -613
rect -119 -629 -41 -613
rect 41 -629 119 -613
rect 201 -629 279 -613
rect -263 -645 -247 -629
rect -233 -645 -217 -629
rect -103 -645 -87 -629
rect -73 -645 -57 -629
rect 57 -645 73 -629
rect 87 -645 103 -629
rect 217 -645 233 -629
rect 247 -645 263 -629
rect -263 -703 -247 -687
rect -233 -703 -217 -687
rect -103 -703 -87 -687
rect -73 -703 -57 -687
rect 57 -703 73 -687
rect 87 -703 103 -687
rect 217 -703 233 -687
rect 247 -703 263 -687
rect -279 -719 -201 -703
rect -119 -719 -41 -703
rect 41 -719 119 -703
rect 201 -719 279 -703
rect -274 -733 -206 -719
rect -114 -733 -46 -719
rect 46 -733 114 -719
rect 206 -733 274 -719
rect -279 -749 -201 -733
rect -119 -749 -41 -733
rect 41 -749 119 -733
rect 201 -749 279 -733
rect -263 -765 -247 -749
rect -233 -765 -217 -749
rect -103 -765 -87 -749
rect -73 -765 -57 -749
rect 57 -765 73 -749
rect 87 -765 103 -749
rect 217 -765 233 -749
rect 247 -765 263 -749
rect -343 -795 -327 -779
rect -313 -795 -297 -779
rect -183 -795 -167 -779
rect -153 -795 -137 -779
rect -23 -795 -7 -779
rect 7 -795 23 -779
rect 137 -795 153 -779
rect 167 -795 183 -779
rect 297 -795 313 -779
rect 327 -795 343 -779
rect -359 -811 -343 -795
rect -297 -811 -281 -795
rect -199 -811 -183 -795
rect -137 -811 -121 -795
rect -39 -811 -23 -795
rect 23 -811 39 -795
rect 121 -811 137 -795
rect 183 -811 199 -795
rect 281 -811 297 -795
rect 343 -811 359 -795
rect -359 -1869 -343 -1853
rect -297 -1868 -281 -1853
rect -199 -1868 -183 -1853
rect -297 -1869 -183 -1868
rect -137 -1868 -121 -1853
rect -39 -1868 -23 -1853
rect -137 -1869 -23 -1868
rect 23 -1868 39 -1853
rect 121 -1868 137 -1853
rect 23 -1869 137 -1868
rect 183 -1868 199 -1853
rect 281 -1868 297 -1853
rect 183 -1869 297 -1868
rect 343 -1869 359 -1853
rect -343 -1885 -327 -1869
rect -313 -1882 -167 -1869
rect -313 -1885 -297 -1882
rect -183 -1885 -167 -1882
rect -153 -1882 -7 -1869
rect -153 -1885 -137 -1882
rect -23 -1885 -7 -1882
rect 7 -1882 153 -1869
rect 7 -1885 23 -1882
rect 137 -1885 153 -1882
rect 167 -1882 313 -1869
rect 167 -1885 183 -1882
rect 297 -1885 313 -1882
rect 327 -1885 343 -1869
rect -263 -1915 -247 -1899
rect -233 -1915 -217 -1899
rect -103 -1915 -87 -1899
rect -73 -1915 -57 -1899
rect 57 -1915 73 -1899
rect 87 -1915 103 -1899
rect 217 -1915 233 -1899
rect 247 -1915 263 -1899
rect -279 -1931 -201 -1915
rect -119 -1931 -41 -1915
rect 41 -1931 119 -1915
rect 201 -1931 279 -1915
rect -274 -1945 -206 -1931
rect -114 -1945 -46 -1931
rect 46 -1945 114 -1931
rect 206 -1945 274 -1931
rect -279 -1961 -201 -1945
rect -119 -1961 -41 -1945
rect 41 -1961 119 -1945
rect 201 -1961 279 -1945
rect -263 -1977 -247 -1961
rect -233 -1977 -217 -1961
rect -103 -1977 -87 -1961
rect -73 -1977 -57 -1961
rect 57 -1977 73 -1961
rect 87 -1977 103 -1961
rect 217 -1977 233 -1961
rect 247 -1977 263 -1961
rect -263 -2035 -247 -2019
rect -233 -2035 -217 -2019
rect -103 -2035 -87 -2019
rect -73 -2035 -57 -2019
rect 57 -2035 73 -2019
rect 87 -2035 103 -2019
rect 217 -2035 233 -2019
rect 247 -2035 263 -2019
rect -279 -2051 -201 -2035
rect -119 -2051 -41 -2035
rect 41 -2051 119 -2035
rect 201 -2051 279 -2035
rect -274 -2065 -206 -2051
rect -114 -2065 -46 -2051
rect 46 -2065 114 -2051
rect 206 -2065 274 -2051
rect -279 -2081 -201 -2065
rect -119 -2081 -41 -2065
rect 41 -2081 119 -2065
rect 201 -2081 279 -2065
rect -263 -2097 -247 -2081
rect -233 -2097 -217 -2081
rect -103 -2097 -87 -2081
rect -73 -2097 -57 -2081
rect 57 -2097 73 -2081
rect 87 -2097 103 -2081
rect 217 -2097 233 -2081
rect 247 -2097 263 -2081
rect -343 -2127 -327 -2111
rect -313 -2127 -297 -2111
rect -183 -2127 -167 -2111
rect -153 -2127 -137 -2111
rect -23 -2127 -7 -2111
rect 7 -2127 23 -2111
rect 137 -2127 153 -2111
rect 167 -2127 183 -2111
rect 297 -2127 313 -2111
rect 327 -2127 343 -2111
rect -359 -2143 -343 -2127
rect -297 -2143 -281 -2127
rect -199 -2143 -183 -2127
rect -137 -2143 -121 -2127
rect -39 -2143 -23 -2127
rect 23 -2143 39 -2127
rect 121 -2143 137 -2127
rect 183 -2143 199 -2127
rect 281 -2143 297 -2127
rect 343 -2143 359 -2127
rect -359 -3201 -343 -3185
rect -297 -3200 -281 -3185
rect -199 -3200 -183 -3185
rect -297 -3201 -183 -3200
rect -137 -3200 -121 -3185
rect -39 -3200 -23 -3185
rect -137 -3201 -23 -3200
rect 23 -3200 39 -3185
rect 121 -3200 137 -3185
rect 23 -3201 137 -3200
rect 183 -3200 199 -3185
rect 281 -3200 297 -3185
rect 183 -3201 297 -3200
rect 343 -3201 359 -3185
rect -343 -3217 -327 -3201
rect -313 -3214 -167 -3201
rect -313 -3217 -297 -3214
rect -183 -3217 -167 -3214
rect -153 -3214 -7 -3201
rect -153 -3217 -137 -3214
rect -23 -3217 -7 -3214
rect 7 -3214 153 -3201
rect 7 -3217 23 -3214
rect 137 -3217 153 -3214
rect 167 -3214 313 -3201
rect 167 -3217 183 -3214
rect 297 -3217 313 -3214
rect 327 -3217 343 -3201
rect -263 -3247 -247 -3231
rect -233 -3247 -217 -3231
rect -103 -3247 -87 -3231
rect -73 -3247 -57 -3231
rect 57 -3247 73 -3231
rect 87 -3247 103 -3231
rect 217 -3247 233 -3231
rect 247 -3247 263 -3231
rect -279 -3263 -201 -3247
rect -119 -3263 -41 -3247
rect 41 -3263 119 -3247
rect 201 -3263 279 -3247
rect -497 -3284 -481 -3268
rect -435 -3284 -419 -3268
rect -274 -3277 -206 -3263
rect -114 -3277 -46 -3263
rect 46 -3277 114 -3263
rect 206 -3277 274 -3263
rect 482 -3268 494 3268
rect -494 -3388 -482 -3284
rect -481 -3300 -465 -3284
rect -451 -3300 -435 -3284
rect -279 -3293 -201 -3277
rect -119 -3293 -41 -3277
rect 41 -3293 119 -3277
rect 201 -3293 279 -3277
rect 419 -3284 435 -3268
rect 481 -3284 497 -3268
rect -263 -3309 -247 -3293
rect -233 -3309 -217 -3293
rect -103 -3309 -87 -3293
rect -73 -3309 -57 -3293
rect 57 -3309 73 -3293
rect 87 -3309 103 -3293
rect 217 -3309 233 -3293
rect 247 -3309 263 -3293
rect 435 -3300 451 -3284
rect 465 -3300 481 -3284
rect 482 -3388 494 -3284
rect -494 -3400 494 -3388
rect 518 -3424 530 3424
rect -530 -3436 530 -3424
<< nwell >>
rect -518 -3424 518 3424
<< pmos >>
rect -268 2114 -212 3214
rect -108 2114 -52 3214
rect 52 2114 108 3214
rect 212 2114 268 3214
rect -268 782 -212 1882
rect -108 782 -52 1882
rect 52 782 108 1882
rect 212 782 268 1882
rect -268 -550 -212 550
rect -108 -550 -52 550
rect 52 -550 108 550
rect 212 -550 268 550
rect -268 -1882 -212 -782
rect -108 -1882 -52 -782
rect 52 -1882 108 -782
rect 212 -1882 268 -782
rect -268 -3214 -212 -2114
rect -108 -3214 -52 -2114
rect 52 -3214 108 -2114
rect 212 -3214 268 -2114
<< pdiff >>
rect -356 3201 -268 3214
rect -356 2127 -343 3201
rect -297 2127 -268 3201
rect -356 2114 -268 2127
rect -212 3201 -108 3214
rect -212 2127 -183 3201
rect -137 2127 -108 3201
rect -212 2114 -108 2127
rect -52 3201 52 3214
rect -52 2127 -23 3201
rect 23 2127 52 3201
rect -52 2114 52 2127
rect 108 3201 212 3214
rect 108 2127 137 3201
rect 183 2127 212 3201
rect 108 2114 212 2127
rect 268 3201 356 3214
rect 268 2127 297 3201
rect 343 2127 356 3201
rect 268 2114 356 2127
rect -356 1869 -268 1882
rect -356 795 -343 1869
rect -297 795 -268 1869
rect -356 782 -268 795
rect -212 1869 -108 1882
rect -212 795 -183 1869
rect -137 795 -108 1869
rect -212 782 -108 795
rect -52 1869 52 1882
rect -52 795 -23 1869
rect 23 795 52 1869
rect -52 782 52 795
rect 108 1869 212 1882
rect 108 795 137 1869
rect 183 795 212 1869
rect 108 782 212 795
rect 268 1869 356 1882
rect 268 795 297 1869
rect 343 795 356 1869
rect 268 782 356 795
rect -356 537 -268 550
rect -356 -537 -343 537
rect -297 -537 -268 537
rect -356 -550 -268 -537
rect -212 537 -108 550
rect -212 -537 -183 537
rect -137 -537 -108 537
rect -212 -550 -108 -537
rect -52 537 52 550
rect -52 -537 -23 537
rect 23 -537 52 537
rect -52 -550 52 -537
rect 108 537 212 550
rect 108 -537 137 537
rect 183 -537 212 537
rect 108 -550 212 -537
rect 268 537 356 550
rect 268 -537 297 537
rect 343 -537 356 537
rect 268 -550 356 -537
rect -356 -795 -268 -782
rect -356 -1869 -343 -795
rect -297 -1869 -268 -795
rect -356 -1882 -268 -1869
rect -212 -795 -108 -782
rect -212 -1869 -183 -795
rect -137 -1869 -108 -795
rect -212 -1882 -108 -1869
rect -52 -795 52 -782
rect -52 -1869 -23 -795
rect 23 -1869 52 -795
rect -52 -1882 52 -1869
rect 108 -795 212 -782
rect 108 -1869 137 -795
rect 183 -1869 212 -795
rect 108 -1882 212 -1869
rect 268 -795 356 -782
rect 268 -1869 297 -795
rect 343 -1869 356 -795
rect 268 -1882 356 -1869
rect -356 -2127 -268 -2114
rect -356 -3201 -343 -2127
rect -297 -3201 -268 -2127
rect -356 -3214 -268 -3201
rect -212 -2127 -108 -2114
rect -212 -3201 -183 -2127
rect -137 -3201 -108 -2127
rect -212 -3214 -108 -3201
rect -52 -2127 52 -2114
rect -52 -3201 -23 -2127
rect 23 -3201 52 -2127
rect -52 -3214 52 -3201
rect 108 -2127 212 -2114
rect 108 -3201 137 -2127
rect 183 -3201 212 -2127
rect 108 -3214 212 -3201
rect 268 -2127 356 -2114
rect 268 -3201 297 -2127
rect 343 -3201 356 -2127
rect 268 -3214 356 -3201
<< pdiffc >>
rect -343 2127 -297 3201
rect -183 2127 -137 3201
rect -23 2127 23 3201
rect 137 2127 183 3201
rect 297 2127 343 3201
rect -343 795 -297 1869
rect -183 795 -137 1869
rect -23 795 23 1869
rect 137 795 183 1869
rect 297 795 343 1869
rect -343 -537 -297 537
rect -183 -537 -137 537
rect -23 -537 23 537
rect 137 -537 183 537
rect 297 -537 343 537
rect -343 -1869 -297 -795
rect -183 -1869 -137 -795
rect -23 -1869 23 -795
rect 137 -1869 183 -795
rect 297 -1869 343 -795
rect -343 -3201 -297 -2127
rect -183 -3201 -137 -2127
rect -23 -3201 23 -2127
rect 137 -3201 183 -2127
rect 297 -3201 343 -2127
<< nsubdiff >>
rect -494 3328 494 3400
rect -494 3284 -422 3328
rect -494 -3284 -481 3284
rect -435 -3284 -422 3284
rect 422 3284 494 3328
rect -494 -3328 -422 -3284
rect 422 -3284 435 3284
rect 481 -3284 494 3284
rect 422 -3328 494 -3284
rect -494 -3400 494 -3328
<< nsubdiffcont >>
rect -481 -3284 -435 3284
rect 435 -3284 481 3284
<< poly >>
rect -276 3293 -204 3306
rect -276 3247 -263 3293
rect -217 3247 -204 3293
rect -276 3234 -204 3247
rect -116 3293 -44 3306
rect -116 3247 -103 3293
rect -57 3247 -44 3293
rect -116 3234 -44 3247
rect 44 3293 116 3306
rect 44 3247 57 3293
rect 103 3247 116 3293
rect 44 3234 116 3247
rect 204 3293 276 3306
rect 204 3247 217 3293
rect 263 3247 276 3293
rect 204 3234 276 3247
rect -268 3214 -212 3234
rect -108 3214 -52 3234
rect 52 3214 108 3234
rect 212 3214 268 3234
rect -268 2094 -212 2114
rect -108 2094 -52 2114
rect 52 2094 108 2114
rect 212 2094 268 2114
rect -276 2081 -204 2094
rect -276 2035 -263 2081
rect -217 2035 -204 2081
rect -276 2022 -204 2035
rect -116 2081 -44 2094
rect -116 2035 -103 2081
rect -57 2035 -44 2081
rect -116 2022 -44 2035
rect 44 2081 116 2094
rect 44 2035 57 2081
rect 103 2035 116 2081
rect 44 2022 116 2035
rect 204 2081 276 2094
rect 204 2035 217 2081
rect 263 2035 276 2081
rect 204 2022 276 2035
rect -276 1961 -204 1974
rect -276 1915 -263 1961
rect -217 1915 -204 1961
rect -276 1902 -204 1915
rect -116 1961 -44 1974
rect -116 1915 -103 1961
rect -57 1915 -44 1961
rect -116 1902 -44 1915
rect 44 1961 116 1974
rect 44 1915 57 1961
rect 103 1915 116 1961
rect 44 1902 116 1915
rect 204 1961 276 1974
rect 204 1915 217 1961
rect 263 1915 276 1961
rect 204 1902 276 1915
rect -268 1882 -212 1902
rect -108 1882 -52 1902
rect 52 1882 108 1902
rect 212 1882 268 1902
rect -268 762 -212 782
rect -108 762 -52 782
rect 52 762 108 782
rect 212 762 268 782
rect -276 749 -204 762
rect -276 703 -263 749
rect -217 703 -204 749
rect -276 690 -204 703
rect -116 749 -44 762
rect -116 703 -103 749
rect -57 703 -44 749
rect -116 690 -44 703
rect 44 749 116 762
rect 44 703 57 749
rect 103 703 116 749
rect 44 690 116 703
rect 204 749 276 762
rect 204 703 217 749
rect 263 703 276 749
rect 204 690 276 703
rect -276 629 -204 642
rect -276 583 -263 629
rect -217 583 -204 629
rect -276 570 -204 583
rect -116 629 -44 642
rect -116 583 -103 629
rect -57 583 -44 629
rect -116 570 -44 583
rect 44 629 116 642
rect 44 583 57 629
rect 103 583 116 629
rect 44 570 116 583
rect 204 629 276 642
rect 204 583 217 629
rect 263 583 276 629
rect 204 570 276 583
rect -268 550 -212 570
rect -108 550 -52 570
rect 52 550 108 570
rect 212 550 268 570
rect -268 -570 -212 -550
rect -108 -570 -52 -550
rect 52 -570 108 -550
rect 212 -570 268 -550
rect -276 -583 -204 -570
rect -276 -629 -263 -583
rect -217 -629 -204 -583
rect -276 -642 -204 -629
rect -116 -583 -44 -570
rect -116 -629 -103 -583
rect -57 -629 -44 -583
rect -116 -642 -44 -629
rect 44 -583 116 -570
rect 44 -629 57 -583
rect 103 -629 116 -583
rect 44 -642 116 -629
rect 204 -583 276 -570
rect 204 -629 217 -583
rect 263 -629 276 -583
rect 204 -642 276 -629
rect -276 -703 -204 -690
rect -276 -749 -263 -703
rect -217 -749 -204 -703
rect -276 -762 -204 -749
rect -116 -703 -44 -690
rect -116 -749 -103 -703
rect -57 -749 -44 -703
rect -116 -762 -44 -749
rect 44 -703 116 -690
rect 44 -749 57 -703
rect 103 -749 116 -703
rect 44 -762 116 -749
rect 204 -703 276 -690
rect 204 -749 217 -703
rect 263 -749 276 -703
rect 204 -762 276 -749
rect -268 -782 -212 -762
rect -108 -782 -52 -762
rect 52 -782 108 -762
rect 212 -782 268 -762
rect -268 -1902 -212 -1882
rect -108 -1902 -52 -1882
rect 52 -1902 108 -1882
rect 212 -1902 268 -1882
rect -276 -1915 -204 -1902
rect -276 -1961 -263 -1915
rect -217 -1961 -204 -1915
rect -276 -1974 -204 -1961
rect -116 -1915 -44 -1902
rect -116 -1961 -103 -1915
rect -57 -1961 -44 -1915
rect -116 -1974 -44 -1961
rect 44 -1915 116 -1902
rect 44 -1961 57 -1915
rect 103 -1961 116 -1915
rect 44 -1974 116 -1961
rect 204 -1915 276 -1902
rect 204 -1961 217 -1915
rect 263 -1961 276 -1915
rect 204 -1974 276 -1961
rect -276 -2035 -204 -2022
rect -276 -2081 -263 -2035
rect -217 -2081 -204 -2035
rect -276 -2094 -204 -2081
rect -116 -2035 -44 -2022
rect -116 -2081 -103 -2035
rect -57 -2081 -44 -2035
rect -116 -2094 -44 -2081
rect 44 -2035 116 -2022
rect 44 -2081 57 -2035
rect 103 -2081 116 -2035
rect 44 -2094 116 -2081
rect 204 -2035 276 -2022
rect 204 -2081 217 -2035
rect 263 -2081 276 -2035
rect 204 -2094 276 -2081
rect -268 -2114 -212 -2094
rect -108 -2114 -52 -2094
rect 52 -2114 108 -2094
rect 212 -2114 268 -2094
rect -268 -3234 -212 -3214
rect -108 -3234 -52 -3214
rect 52 -3234 108 -3214
rect 212 -3234 268 -3214
rect -276 -3247 -204 -3234
rect -276 -3293 -263 -3247
rect -217 -3293 -204 -3247
rect -276 -3306 -204 -3293
rect -116 -3247 -44 -3234
rect -116 -3293 -103 -3247
rect -57 -3293 -44 -3247
rect -116 -3306 -44 -3293
rect 44 -3247 116 -3234
rect 44 -3293 57 -3247
rect 103 -3293 116 -3247
rect 44 -3306 116 -3293
rect 204 -3247 276 -3234
rect 204 -3293 217 -3247
rect 263 -3293 276 -3247
rect 204 -3306 276 -3293
<< polycont >>
rect -263 3247 -217 3293
rect -103 3247 -57 3293
rect 57 3247 103 3293
rect 217 3247 263 3293
rect -263 2035 -217 2081
rect -103 2035 -57 2081
rect 57 2035 103 2081
rect 217 2035 263 2081
rect -263 1915 -217 1961
rect -103 1915 -57 1961
rect 57 1915 103 1961
rect 217 1915 263 1961
rect -263 703 -217 749
rect -103 703 -57 749
rect 57 703 103 749
rect 217 703 263 749
rect -263 583 -217 629
rect -103 583 -57 629
rect 57 583 103 629
rect 217 583 263 629
rect -263 -629 -217 -583
rect -103 -629 -57 -583
rect 57 -629 103 -583
rect 217 -629 263 -583
rect -263 -749 -217 -703
rect -103 -749 -57 -703
rect 57 -749 103 -703
rect 217 -749 263 -703
rect -263 -1961 -217 -1915
rect -103 -1961 -57 -1915
rect 57 -1961 103 -1915
rect 217 -1961 263 -1915
rect -263 -2081 -217 -2035
rect -103 -2081 -57 -2035
rect 57 -2081 103 -2035
rect 217 -2081 263 -2035
rect -263 -3293 -217 -3247
rect -103 -3293 -57 -3247
rect 57 -3293 103 -3247
rect 217 -3293 263 -3247
<< metal1 >>
rect -481 3341 481 3387
rect -481 -3341 -435 3341
rect -274 3247 -206 3293
rect -114 3247 -46 3293
rect 46 3247 114 3293
rect 206 3247 274 3293
rect -343 2116 -297 3212
rect -183 2116 -137 3212
rect -23 2116 23 3212
rect 137 2116 183 3212
rect 297 2116 343 3212
rect -274 2035 -206 2081
rect -114 2035 -46 2081
rect 46 2035 114 2081
rect 206 2035 274 2081
rect -274 1915 -206 1961
rect -114 1915 -46 1961
rect 46 1915 114 1961
rect 206 1915 274 1961
rect -343 784 -297 1880
rect -183 784 -137 1880
rect -23 784 23 1880
rect 137 784 183 1880
rect 297 784 343 1880
rect -274 703 -206 749
rect -114 703 -46 749
rect 46 703 114 749
rect 206 703 274 749
rect -274 583 -206 629
rect -114 583 -46 629
rect 46 583 114 629
rect 206 583 274 629
rect -343 -548 -297 548
rect -183 -548 -137 548
rect -23 -548 23 548
rect 137 -548 183 548
rect 297 -548 343 548
rect -274 -629 -206 -583
rect -114 -629 -46 -583
rect 46 -629 114 -583
rect 206 -629 274 -583
rect -274 -749 -206 -703
rect -114 -749 -46 -703
rect 46 -749 114 -703
rect 206 -749 274 -703
rect -343 -1880 -297 -784
rect -183 -1880 -137 -784
rect -23 -1880 23 -784
rect 137 -1880 183 -784
rect 297 -1880 343 -784
rect -274 -1961 -206 -1915
rect -114 -1961 -46 -1915
rect 46 -1961 114 -1915
rect 206 -1961 274 -1915
rect -274 -2081 -206 -2035
rect -114 -2081 -46 -2035
rect 46 -2081 114 -2035
rect 206 -2081 274 -2035
rect -343 -3212 -297 -2116
rect -183 -3212 -137 -2116
rect -23 -3212 23 -2116
rect 137 -3212 183 -2116
rect 297 -3212 343 -2116
rect -274 -3293 -206 -3247
rect -114 -3293 -46 -3247
rect 46 -3293 114 -3247
rect 206 -3293 274 -3247
rect 435 -3341 481 3341
rect -481 -3387 481 -3341
<< properties >>
string FIXED_BBOX -458 -3364 458 3364
string gencell pfet_03v3
string library gf180mcu
string parameters w 5.5 l 0.280 m 5 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 class mosfet full_metal 1 compatible {pfet_03v3 pfet_06v0}
<< end >>

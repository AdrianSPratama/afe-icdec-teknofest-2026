magic
tech sky130A
magscale 1 2
timestamp 1771462974
<< error_p >>
rect -29 166 29 172
rect -29 132 -17 166
rect -29 126 29 132
<< nmos >>
rect -30 -156 30 94
<< ndiff >>
rect -88 82 -30 94
rect -88 -144 -76 82
rect -42 -144 -30 82
rect -88 -156 -30 -144
rect 30 82 88 94
rect 30 -144 42 82
rect 76 -144 88 82
rect 30 -156 88 -144
<< ndiffc >>
rect -76 -144 -42 82
rect 42 -144 76 82
<< poly >>
rect -33 166 33 182
rect -33 132 -17 166
rect 17 132 33 166
rect -33 116 33 132
rect -30 94 30 116
rect -30 -182 30 -156
<< polycont >>
rect -17 132 17 166
<< locali >>
rect -33 132 -17 166
rect 17 132 33 166
rect -76 82 -42 98
rect -76 -160 -42 -144
rect 42 82 76 98
rect 42 -160 76 -144
<< viali >>
rect -17 132 17 166
rect -76 -144 -42 82
rect 42 -144 76 82
<< metal1 >>
rect -29 166 29 172
rect -29 132 -17 166
rect 17 132 29 166
rect -29 126 29 132
rect -82 82 -36 94
rect -82 -144 -76 82
rect -42 -144 -36 82
rect -82 -156 -36 -144
rect 36 82 82 94
rect 36 -144 42 82
rect 76 -144 82 82
rect 36 -156 82 -144
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1.25 l 0.3 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 class mosfet compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

** sch_path: /foss/designs/afe-icdec-teknofest-2026/bandgap/bgr/current-mode-bgr.sch
.subckt current-mode-bgr IREF VDD VSS
*.PININFO IREF:O VDD:B VSS:B
R21 VSS net1 sky130_fd_pr__res_generic_l1 W=1 L=4.1 m=1
R1 VSS net1 sky130_fd_pr__res_generic_l1 W=1 L=4.1 m=1
R3 VSS net1 sky130_fd_pr__res_generic_l1 W=1 L=4.1 m=1
R4 VSS net1 sky130_fd_pr__res_generic_l1 W=1 L=4.1 m=1
R5 VSS net1 sky130_fd_pr__res_generic_l1 W=1 L=4.1 m=1
R6 VSS net1 sky130_fd_pr__res_generic_l1 W=1 L=4.1 m=1
R7 VSS net1 sky130_fd_pr__res_generic_l1 W=1 L=4.1 m=1
R8 VSS net1 sky130_fd_pr__res_generic_l1 W=1 L=4.1 m=1
R9 VSS net1 sky130_fd_pr__res_generic_l1 W=1 L=4.1 m=1
R10 VSS net1 sky130_fd_pr__res_generic_l1 W=1 L=4.1 m=1
XR11 net3 net2 VSS sky130_fd_pr__res_xhigh_po_1p41 L=1.41 mult=1 m=1
XR2 net5 net3 VSS sky130_fd_pr__res_xhigh_po_1p41 L=1.41 mult=1 m=1
XR12 net4 net5 VSS sky130_fd_pr__res_xhigh_po_1p41 L=1.41 mult=1 m=1
XR13 net11 net4 VSS sky130_fd_pr__res_xhigh_po_1p41 L=1.41 mult=1 m=1
XR14 net6 net11 VSS sky130_fd_pr__res_xhigh_po_1p41 L=1.41 mult=1 m=1
XR15 net10 net6 VSS sky130_fd_pr__res_xhigh_po_1p41 L=1.41 mult=1 m=1
XR16 net7 net10 VSS sky130_fd_pr__res_xhigh_po_1p41 L=1.41 mult=1 m=1
XR17 net9 net7 VSS sky130_fd_pr__res_xhigh_po_1p41 L=1.41 mult=1 m=1
XR18 net8 net9 VSS sky130_fd_pr__res_xhigh_po_1p41 L=1.41 mult=1 m=1
XR19 VSS net8 VSS sky130_fd_pr__res_xhigh_po_1p41 L=1.41 mult=1 m=1
XM14 net12 net13 net1 VSS sky130_fd_pr__nfet_01v8 L=5 W=10 nf=4 m=1
XM15 net13 net13 VSS VSS sky130_fd_pr__nfet_01v8 L=5 W=10 nf=4 m=1
XM16 net12 net12 VDD VDD sky130_fd_pr__pfet_01v8 L=5 W=20 nf=2 m=1
XM17 net13 net12 VDD VDD sky130_fd_pr__pfet_01v8 L=5 W=20 nf=2 m=1
XM18 net13 VSS VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 m=1
XM19 VSS net12 VDD VDD sky130_fd_pr__pfet_01v8 L=1.5 W=20 nf=4 m=1
XM20 VSS net12 VDD VDD sky130_fd_pr__pfet_01v8 L=1.5 W=20 nf=4 m=1
XM21 net14 net14 VDD VDD sky130_fd_pr__pfet_01v8 L=1.5 W=2 nf=1 m=1
XM22 net2 net14 VDD VDD sky130_fd_pr__pfet_01v8 L=1.5 W=2 nf=1 m=1
XM23 IREF net12 VDD VDD sky130_fd_pr__pfet_01v8 L=5 W=6.35 nf=1 m=1
XM24 IREF net14 VDD VDD sky130_fd_pr__pfet_01v8 L=5 W=25 nf=4 m=1
XM25 net14 VSS VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XM26 VSS net2 VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
.ends

magic
tech sky130A
magscale 1 2
timestamp 1771413069
<< error_p >>
rect -681 2022 681 2240
rect -681 686 681 904
rect -681 -650 681 -432
rect -681 -1986 681 -1768
<< nwell >>
rect -681 2022 681 3322
rect -681 686 681 1986
rect -681 -650 681 650
rect -681 -1986 681 -686
rect -681 -3322 681 -2022
<< pmos >>
rect -587 2122 -337 3222
rect -279 2122 -29 3222
rect 29 2122 279 3222
rect 337 2122 587 3222
rect -587 786 -337 1886
rect -279 786 -29 1886
rect 29 786 279 1886
rect 337 786 587 1886
rect -587 -550 -337 550
rect -279 -550 -29 550
rect 29 -550 279 550
rect 337 -550 587 550
rect -587 -1886 -337 -786
rect -279 -1886 -29 -786
rect 29 -1886 279 -786
rect 337 -1886 587 -786
rect -587 -3222 -337 -2122
rect -279 -3222 -29 -2122
rect 29 -3222 279 -2122
rect 337 -3222 587 -2122
<< pdiff >>
rect -645 3210 -587 3222
rect -645 2134 -633 3210
rect -599 2134 -587 3210
rect -645 2122 -587 2134
rect -337 3210 -279 3222
rect -337 2134 -325 3210
rect -291 2134 -279 3210
rect -337 2122 -279 2134
rect -29 3210 29 3222
rect -29 2134 -17 3210
rect 17 2134 29 3210
rect -29 2122 29 2134
rect 279 3210 337 3222
rect 279 2134 291 3210
rect 325 2134 337 3210
rect 279 2122 337 2134
rect 587 3210 645 3222
rect 587 2134 599 3210
rect 633 2134 645 3210
rect 587 2122 645 2134
rect -645 1874 -587 1886
rect -645 798 -633 1874
rect -599 798 -587 1874
rect -645 786 -587 798
rect -337 1874 -279 1886
rect -337 798 -325 1874
rect -291 798 -279 1874
rect -337 786 -279 798
rect -29 1874 29 1886
rect -29 798 -17 1874
rect 17 798 29 1874
rect -29 786 29 798
rect 279 1874 337 1886
rect 279 798 291 1874
rect 325 798 337 1874
rect 279 786 337 798
rect 587 1874 645 1886
rect 587 798 599 1874
rect 633 798 645 1874
rect 587 786 645 798
rect -645 538 -587 550
rect -645 -538 -633 538
rect -599 -538 -587 538
rect -645 -550 -587 -538
rect -337 538 -279 550
rect -337 -538 -325 538
rect -291 -538 -279 538
rect -337 -550 -279 -538
rect -29 538 29 550
rect -29 -538 -17 538
rect 17 -538 29 538
rect -29 -550 29 -538
rect 279 538 337 550
rect 279 -538 291 538
rect 325 -538 337 538
rect 279 -550 337 -538
rect 587 538 645 550
rect 587 -538 599 538
rect 633 -538 645 538
rect 587 -550 645 -538
rect -645 -798 -587 -786
rect -645 -1874 -633 -798
rect -599 -1874 -587 -798
rect -645 -1886 -587 -1874
rect -337 -798 -279 -786
rect -337 -1874 -325 -798
rect -291 -1874 -279 -798
rect -337 -1886 -279 -1874
rect -29 -798 29 -786
rect -29 -1874 -17 -798
rect 17 -1874 29 -798
rect -29 -1886 29 -1874
rect 279 -798 337 -786
rect 279 -1874 291 -798
rect 325 -1874 337 -798
rect 279 -1886 337 -1874
rect 587 -798 645 -786
rect 587 -1874 599 -798
rect 633 -1874 645 -798
rect 587 -1886 645 -1874
rect -645 -2134 -587 -2122
rect -645 -3210 -633 -2134
rect -599 -3210 -587 -2134
rect -645 -3222 -587 -3210
rect -337 -2134 -279 -2122
rect -337 -3210 -325 -2134
rect -291 -3210 -279 -2134
rect -337 -3222 -279 -3210
rect -29 -2134 29 -2122
rect -29 -3210 -17 -2134
rect 17 -3210 29 -2134
rect -29 -3222 29 -3210
rect 279 -2134 337 -2122
rect 279 -3210 291 -2134
rect 325 -3210 337 -2134
rect 279 -3222 337 -3210
rect 587 -2134 645 -2122
rect 587 -3210 599 -2134
rect 633 -3210 645 -2134
rect 587 -3222 645 -3210
<< pdiffc >>
rect -633 2134 -599 3210
rect -325 2134 -291 3210
rect -17 2134 17 3210
rect 291 2134 325 3210
rect 599 2134 633 3210
rect -633 798 -599 1874
rect -325 798 -291 1874
rect -17 798 17 1874
rect 291 798 325 1874
rect 599 798 633 1874
rect -633 -538 -599 538
rect -325 -538 -291 538
rect -17 -538 17 538
rect 291 -538 325 538
rect 599 -538 633 538
rect -633 -1874 -599 -798
rect -325 -1874 -291 -798
rect -17 -1874 17 -798
rect 291 -1874 325 -798
rect 599 -1874 633 -798
rect -633 -3210 -599 -2134
rect -325 -3210 -291 -2134
rect -17 -3210 17 -2134
rect 291 -3210 325 -2134
rect 599 -3210 633 -2134
<< poly >>
rect -587 3303 -337 3319
rect -587 3269 -571 3303
rect -353 3269 -337 3303
rect -587 3222 -337 3269
rect -279 3303 -29 3319
rect -279 3269 -263 3303
rect -45 3269 -29 3303
rect -279 3222 -29 3269
rect 29 3303 279 3319
rect 29 3269 45 3303
rect 263 3269 279 3303
rect 29 3222 279 3269
rect 337 3303 587 3319
rect 337 3269 353 3303
rect 571 3269 587 3303
rect 337 3222 587 3269
rect -587 2075 -337 2122
rect -587 2041 -571 2075
rect -353 2041 -337 2075
rect -587 2025 -337 2041
rect -279 2075 -29 2122
rect -279 2041 -263 2075
rect -45 2041 -29 2075
rect -279 2025 -29 2041
rect 29 2075 279 2122
rect 29 2041 45 2075
rect 263 2041 279 2075
rect 29 2025 279 2041
rect 337 2075 587 2122
rect 337 2041 353 2075
rect 571 2041 587 2075
rect 337 2025 587 2041
rect -587 1967 -337 1983
rect -587 1933 -571 1967
rect -353 1933 -337 1967
rect -587 1886 -337 1933
rect -279 1967 -29 1983
rect -279 1933 -263 1967
rect -45 1933 -29 1967
rect -279 1886 -29 1933
rect 29 1967 279 1983
rect 29 1933 45 1967
rect 263 1933 279 1967
rect 29 1886 279 1933
rect 337 1967 587 1983
rect 337 1933 353 1967
rect 571 1933 587 1967
rect 337 1886 587 1933
rect -587 739 -337 786
rect -587 705 -571 739
rect -353 705 -337 739
rect -587 689 -337 705
rect -279 739 -29 786
rect -279 705 -263 739
rect -45 705 -29 739
rect -279 689 -29 705
rect 29 739 279 786
rect 29 705 45 739
rect 263 705 279 739
rect 29 689 279 705
rect 337 739 587 786
rect 337 705 353 739
rect 571 705 587 739
rect 337 689 587 705
rect -587 631 -337 647
rect -587 597 -571 631
rect -353 597 -337 631
rect -587 550 -337 597
rect -279 631 -29 647
rect -279 597 -263 631
rect -45 597 -29 631
rect -279 550 -29 597
rect 29 631 279 647
rect 29 597 45 631
rect 263 597 279 631
rect 29 550 279 597
rect 337 631 587 647
rect 337 597 353 631
rect 571 597 587 631
rect 337 550 587 597
rect -587 -597 -337 -550
rect -587 -631 -571 -597
rect -353 -631 -337 -597
rect -587 -647 -337 -631
rect -279 -597 -29 -550
rect -279 -631 -263 -597
rect -45 -631 -29 -597
rect -279 -647 -29 -631
rect 29 -597 279 -550
rect 29 -631 45 -597
rect 263 -631 279 -597
rect 29 -647 279 -631
rect 337 -597 587 -550
rect 337 -631 353 -597
rect 571 -631 587 -597
rect 337 -647 587 -631
rect -587 -705 -337 -689
rect -587 -739 -571 -705
rect -353 -739 -337 -705
rect -587 -786 -337 -739
rect -279 -705 -29 -689
rect -279 -739 -263 -705
rect -45 -739 -29 -705
rect -279 -786 -29 -739
rect 29 -705 279 -689
rect 29 -739 45 -705
rect 263 -739 279 -705
rect 29 -786 279 -739
rect 337 -705 587 -689
rect 337 -739 353 -705
rect 571 -739 587 -705
rect 337 -786 587 -739
rect -587 -1933 -337 -1886
rect -587 -1967 -571 -1933
rect -353 -1967 -337 -1933
rect -587 -1983 -337 -1967
rect -279 -1933 -29 -1886
rect -279 -1967 -263 -1933
rect -45 -1967 -29 -1933
rect -279 -1983 -29 -1967
rect 29 -1933 279 -1886
rect 29 -1967 45 -1933
rect 263 -1967 279 -1933
rect 29 -1983 279 -1967
rect 337 -1933 587 -1886
rect 337 -1967 353 -1933
rect 571 -1967 587 -1933
rect 337 -1983 587 -1967
rect -587 -2041 -337 -2025
rect -587 -2075 -571 -2041
rect -353 -2075 -337 -2041
rect -587 -2122 -337 -2075
rect -279 -2041 -29 -2025
rect -279 -2075 -263 -2041
rect -45 -2075 -29 -2041
rect -279 -2122 -29 -2075
rect 29 -2041 279 -2025
rect 29 -2075 45 -2041
rect 263 -2075 279 -2041
rect 29 -2122 279 -2075
rect 337 -2041 587 -2025
rect 337 -2075 353 -2041
rect 571 -2075 587 -2041
rect 337 -2122 587 -2075
rect -587 -3269 -337 -3222
rect -587 -3303 -571 -3269
rect -353 -3303 -337 -3269
rect -587 -3319 -337 -3303
rect -279 -3269 -29 -3222
rect -279 -3303 -263 -3269
rect -45 -3303 -29 -3269
rect -279 -3319 -29 -3303
rect 29 -3269 279 -3222
rect 29 -3303 45 -3269
rect 263 -3303 279 -3269
rect 29 -3319 279 -3303
rect 337 -3269 587 -3222
rect 337 -3303 353 -3269
rect 571 -3303 587 -3269
rect 337 -3319 587 -3303
<< polycont >>
rect -571 3269 -353 3303
rect -263 3269 -45 3303
rect 45 3269 263 3303
rect 353 3269 571 3303
rect -571 2041 -353 2075
rect -263 2041 -45 2075
rect 45 2041 263 2075
rect 353 2041 571 2075
rect -571 1933 -353 1967
rect -263 1933 -45 1967
rect 45 1933 263 1967
rect 353 1933 571 1967
rect -571 705 -353 739
rect -263 705 -45 739
rect 45 705 263 739
rect 353 705 571 739
rect -571 597 -353 631
rect -263 597 -45 631
rect 45 597 263 631
rect 353 597 571 631
rect -571 -631 -353 -597
rect -263 -631 -45 -597
rect 45 -631 263 -597
rect 353 -631 571 -597
rect -571 -739 -353 -705
rect -263 -739 -45 -705
rect 45 -739 263 -705
rect 353 -739 571 -705
rect -571 -1967 -353 -1933
rect -263 -1967 -45 -1933
rect 45 -1967 263 -1933
rect 353 -1967 571 -1933
rect -571 -2075 -353 -2041
rect -263 -2075 -45 -2041
rect 45 -2075 263 -2041
rect 353 -2075 571 -2041
rect -571 -3303 -353 -3269
rect -263 -3303 -45 -3269
rect 45 -3303 263 -3269
rect 353 -3303 571 -3269
<< locali >>
rect -587 3269 -571 3303
rect -353 3269 -337 3303
rect -279 3269 -263 3303
rect -45 3269 -29 3303
rect 29 3269 45 3303
rect 263 3269 279 3303
rect 337 3269 353 3303
rect 571 3269 587 3303
rect -633 3210 -599 3226
rect -633 2118 -599 2134
rect -325 3210 -291 3226
rect -325 2118 -291 2134
rect -17 3210 17 3226
rect -17 2118 17 2134
rect 291 3210 325 3226
rect 291 2118 325 2134
rect 599 3210 633 3226
rect 599 2118 633 2134
rect -587 2041 -571 2075
rect -353 2041 -337 2075
rect -279 2041 -263 2075
rect -45 2041 -29 2075
rect 29 2041 45 2075
rect 263 2041 279 2075
rect 337 2041 353 2075
rect 571 2041 587 2075
rect -587 1933 -571 1967
rect -353 1933 -337 1967
rect -279 1933 -263 1967
rect -45 1933 -29 1967
rect 29 1933 45 1967
rect 263 1933 279 1967
rect 337 1933 353 1967
rect 571 1933 587 1967
rect -633 1874 -599 1890
rect -633 782 -599 798
rect -325 1874 -291 1890
rect -325 782 -291 798
rect -17 1874 17 1890
rect -17 782 17 798
rect 291 1874 325 1890
rect 291 782 325 798
rect 599 1874 633 1890
rect 599 782 633 798
rect -587 705 -571 739
rect -353 705 -337 739
rect -279 705 -263 739
rect -45 705 -29 739
rect 29 705 45 739
rect 263 705 279 739
rect 337 705 353 739
rect 571 705 587 739
rect -587 597 -571 631
rect -353 597 -337 631
rect -279 597 -263 631
rect -45 597 -29 631
rect 29 597 45 631
rect 263 597 279 631
rect 337 597 353 631
rect 571 597 587 631
rect -633 538 -599 554
rect -633 -554 -599 -538
rect -325 538 -291 554
rect -325 -554 -291 -538
rect -17 538 17 554
rect -17 -554 17 -538
rect 291 538 325 554
rect 291 -554 325 -538
rect 599 538 633 554
rect 599 -554 633 -538
rect -587 -631 -571 -597
rect -353 -631 -337 -597
rect -279 -631 -263 -597
rect -45 -631 -29 -597
rect 29 -631 45 -597
rect 263 -631 279 -597
rect 337 -631 353 -597
rect 571 -631 587 -597
rect -587 -739 -571 -705
rect -353 -739 -337 -705
rect -279 -739 -263 -705
rect -45 -739 -29 -705
rect 29 -739 45 -705
rect 263 -739 279 -705
rect 337 -739 353 -705
rect 571 -739 587 -705
rect -633 -798 -599 -782
rect -633 -1890 -599 -1874
rect -325 -798 -291 -782
rect -325 -1890 -291 -1874
rect -17 -798 17 -782
rect -17 -1890 17 -1874
rect 291 -798 325 -782
rect 291 -1890 325 -1874
rect 599 -798 633 -782
rect 599 -1890 633 -1874
rect -587 -1967 -571 -1933
rect -353 -1967 -337 -1933
rect -279 -1967 -263 -1933
rect -45 -1967 -29 -1933
rect 29 -1967 45 -1933
rect 263 -1967 279 -1933
rect 337 -1967 353 -1933
rect 571 -1967 587 -1933
rect -587 -2075 -571 -2041
rect -353 -2075 -337 -2041
rect -279 -2075 -263 -2041
rect -45 -2075 -29 -2041
rect 29 -2075 45 -2041
rect 263 -2075 279 -2041
rect 337 -2075 353 -2041
rect 571 -2075 587 -2041
rect -633 -2134 -599 -2118
rect -633 -3226 -599 -3210
rect -325 -2134 -291 -2118
rect -325 -3226 -291 -3210
rect -17 -2134 17 -2118
rect -17 -3226 17 -3210
rect 291 -2134 325 -2118
rect 291 -3226 325 -3210
rect 599 -2134 633 -2118
rect 599 -3226 633 -3210
rect -587 -3303 -571 -3269
rect -353 -3303 -337 -3269
rect -279 -3303 -263 -3269
rect -45 -3303 -29 -3269
rect 29 -3303 45 -3269
rect 263 -3303 279 -3269
rect 337 -3303 353 -3269
rect 571 -3303 587 -3269
<< viali >>
rect -571 3269 -353 3303
rect -263 3269 -45 3303
rect 45 3269 263 3303
rect 353 3269 571 3303
rect -633 2134 -599 3210
rect -325 2134 -291 3210
rect -17 2134 17 3210
rect 291 2134 325 3210
rect 599 2134 633 3210
rect -571 2041 -353 2075
rect -263 2041 -45 2075
rect 45 2041 263 2075
rect 353 2041 571 2075
rect -571 1933 -353 1967
rect -263 1933 -45 1967
rect 45 1933 263 1967
rect 353 1933 571 1967
rect -633 798 -599 1874
rect -325 798 -291 1874
rect -17 798 17 1874
rect 291 798 325 1874
rect 599 798 633 1874
rect -571 705 -353 739
rect -263 705 -45 739
rect 45 705 263 739
rect 353 705 571 739
rect -571 597 -353 631
rect -263 597 -45 631
rect 45 597 263 631
rect 353 597 571 631
rect -633 -538 -599 538
rect -325 -538 -291 538
rect -17 -538 17 538
rect 291 -538 325 538
rect 599 -538 633 538
rect -571 -631 -353 -597
rect -263 -631 -45 -597
rect 45 -631 263 -597
rect 353 -631 571 -597
rect -571 -739 -353 -705
rect -263 -739 -45 -705
rect 45 -739 263 -705
rect 353 -739 571 -705
rect -633 -1874 -599 -798
rect -325 -1874 -291 -798
rect -17 -1874 17 -798
rect 291 -1874 325 -798
rect 599 -1874 633 -798
rect -571 -1967 -353 -1933
rect -263 -1967 -45 -1933
rect 45 -1967 263 -1933
rect 353 -1967 571 -1933
rect -571 -2075 -353 -2041
rect -263 -2075 -45 -2041
rect 45 -2075 263 -2041
rect 353 -2075 571 -2041
rect -633 -3210 -599 -2134
rect -325 -3210 -291 -2134
rect -17 -3210 17 -2134
rect 291 -3210 325 -2134
rect 599 -3210 633 -2134
rect -571 -3303 -353 -3269
rect -263 -3303 -45 -3269
rect 45 -3303 263 -3269
rect 353 -3303 571 -3269
<< metal1 >>
rect -583 3303 -341 3309
rect -583 3269 -571 3303
rect -353 3269 -341 3303
rect -583 3263 -341 3269
rect -275 3303 -33 3309
rect -275 3269 -263 3303
rect -45 3269 -33 3303
rect -275 3263 -33 3269
rect 33 3303 275 3309
rect 33 3269 45 3303
rect 263 3269 275 3303
rect 33 3263 275 3269
rect 341 3303 583 3309
rect 341 3269 353 3303
rect 571 3269 583 3303
rect 341 3263 583 3269
rect -639 3210 -593 3222
rect -639 2134 -633 3210
rect -599 2134 -593 3210
rect -639 2122 -593 2134
rect -331 3210 -285 3222
rect -331 2134 -325 3210
rect -291 2134 -285 3210
rect -331 2122 -285 2134
rect -23 3210 23 3222
rect -23 2134 -17 3210
rect 17 2134 23 3210
rect -23 2122 23 2134
rect 285 3210 331 3222
rect 285 2134 291 3210
rect 325 2134 331 3210
rect 285 2122 331 2134
rect 593 3210 639 3222
rect 593 2134 599 3210
rect 633 2134 639 3210
rect 593 2122 639 2134
rect -583 2075 -341 2081
rect -583 2041 -571 2075
rect -353 2041 -341 2075
rect -583 2035 -341 2041
rect -275 2075 -33 2081
rect -275 2041 -263 2075
rect -45 2041 -33 2075
rect -275 2035 -33 2041
rect 33 2075 275 2081
rect 33 2041 45 2075
rect 263 2041 275 2075
rect 33 2035 275 2041
rect 341 2075 583 2081
rect 341 2041 353 2075
rect 571 2041 583 2075
rect 341 2035 583 2041
rect -583 1967 -341 1973
rect -583 1933 -571 1967
rect -353 1933 -341 1967
rect -583 1927 -341 1933
rect -275 1967 -33 1973
rect -275 1933 -263 1967
rect -45 1933 -33 1967
rect -275 1927 -33 1933
rect 33 1967 275 1973
rect 33 1933 45 1967
rect 263 1933 275 1967
rect 33 1927 275 1933
rect 341 1967 583 1973
rect 341 1933 353 1967
rect 571 1933 583 1967
rect 341 1927 583 1933
rect -639 1874 -593 1886
rect -639 798 -633 1874
rect -599 798 -593 1874
rect -639 786 -593 798
rect -331 1874 -285 1886
rect -331 798 -325 1874
rect -291 798 -285 1874
rect -331 786 -285 798
rect -23 1874 23 1886
rect -23 798 -17 1874
rect 17 798 23 1874
rect -23 786 23 798
rect 285 1874 331 1886
rect 285 798 291 1874
rect 325 798 331 1874
rect 285 786 331 798
rect 593 1874 639 1886
rect 593 798 599 1874
rect 633 798 639 1874
rect 593 786 639 798
rect -583 739 -341 745
rect -583 705 -571 739
rect -353 705 -341 739
rect -583 699 -341 705
rect -275 739 -33 745
rect -275 705 -263 739
rect -45 705 -33 739
rect -275 699 -33 705
rect 33 739 275 745
rect 33 705 45 739
rect 263 705 275 739
rect 33 699 275 705
rect 341 739 583 745
rect 341 705 353 739
rect 571 705 583 739
rect 341 699 583 705
rect -583 631 -341 637
rect -583 597 -571 631
rect -353 597 -341 631
rect -583 591 -341 597
rect -275 631 -33 637
rect -275 597 -263 631
rect -45 597 -33 631
rect -275 591 -33 597
rect 33 631 275 637
rect 33 597 45 631
rect 263 597 275 631
rect 33 591 275 597
rect 341 631 583 637
rect 341 597 353 631
rect 571 597 583 631
rect 341 591 583 597
rect -639 538 -593 550
rect -639 -538 -633 538
rect -599 -538 -593 538
rect -639 -550 -593 -538
rect -331 538 -285 550
rect -331 -538 -325 538
rect -291 -538 -285 538
rect -331 -550 -285 -538
rect -23 538 23 550
rect -23 -538 -17 538
rect 17 -538 23 538
rect -23 -550 23 -538
rect 285 538 331 550
rect 285 -538 291 538
rect 325 -538 331 538
rect 285 -550 331 -538
rect 593 538 639 550
rect 593 -538 599 538
rect 633 -538 639 538
rect 593 -550 639 -538
rect -583 -597 -341 -591
rect -583 -631 -571 -597
rect -353 -631 -341 -597
rect -583 -637 -341 -631
rect -275 -597 -33 -591
rect -275 -631 -263 -597
rect -45 -631 -33 -597
rect -275 -637 -33 -631
rect 33 -597 275 -591
rect 33 -631 45 -597
rect 263 -631 275 -597
rect 33 -637 275 -631
rect 341 -597 583 -591
rect 341 -631 353 -597
rect 571 -631 583 -597
rect 341 -637 583 -631
rect -583 -705 -341 -699
rect -583 -739 -571 -705
rect -353 -739 -341 -705
rect -583 -745 -341 -739
rect -275 -705 -33 -699
rect -275 -739 -263 -705
rect -45 -739 -33 -705
rect -275 -745 -33 -739
rect 33 -705 275 -699
rect 33 -739 45 -705
rect 263 -739 275 -705
rect 33 -745 275 -739
rect 341 -705 583 -699
rect 341 -739 353 -705
rect 571 -739 583 -705
rect 341 -745 583 -739
rect -639 -798 -593 -786
rect -639 -1874 -633 -798
rect -599 -1874 -593 -798
rect -639 -1886 -593 -1874
rect -331 -798 -285 -786
rect -331 -1874 -325 -798
rect -291 -1874 -285 -798
rect -331 -1886 -285 -1874
rect -23 -798 23 -786
rect -23 -1874 -17 -798
rect 17 -1874 23 -798
rect -23 -1886 23 -1874
rect 285 -798 331 -786
rect 285 -1874 291 -798
rect 325 -1874 331 -798
rect 285 -1886 331 -1874
rect 593 -798 639 -786
rect 593 -1874 599 -798
rect 633 -1874 639 -798
rect 593 -1886 639 -1874
rect -583 -1933 -341 -1927
rect -583 -1967 -571 -1933
rect -353 -1967 -341 -1933
rect -583 -1973 -341 -1967
rect -275 -1933 -33 -1927
rect -275 -1967 -263 -1933
rect -45 -1967 -33 -1933
rect -275 -1973 -33 -1967
rect 33 -1933 275 -1927
rect 33 -1967 45 -1933
rect 263 -1967 275 -1933
rect 33 -1973 275 -1967
rect 341 -1933 583 -1927
rect 341 -1967 353 -1933
rect 571 -1967 583 -1933
rect 341 -1973 583 -1967
rect -583 -2041 -341 -2035
rect -583 -2075 -571 -2041
rect -353 -2075 -341 -2041
rect -583 -2081 -341 -2075
rect -275 -2041 -33 -2035
rect -275 -2075 -263 -2041
rect -45 -2075 -33 -2041
rect -275 -2081 -33 -2075
rect 33 -2041 275 -2035
rect 33 -2075 45 -2041
rect 263 -2075 275 -2041
rect 33 -2081 275 -2075
rect 341 -2041 583 -2035
rect 341 -2075 353 -2041
rect 571 -2075 583 -2041
rect 341 -2081 583 -2075
rect -639 -2134 -593 -2122
rect -639 -3210 -633 -2134
rect -599 -3210 -593 -2134
rect -639 -3222 -593 -3210
rect -331 -2134 -285 -2122
rect -331 -3210 -325 -2134
rect -291 -3210 -285 -2134
rect -331 -3222 -285 -3210
rect -23 -2134 23 -2122
rect -23 -3210 -17 -2134
rect 17 -3210 23 -2134
rect -23 -3222 23 -3210
rect 285 -2134 331 -2122
rect 285 -3210 291 -2134
rect 325 -3210 331 -2134
rect 285 -3222 331 -3210
rect 593 -2134 639 -2122
rect 593 -3210 599 -2134
rect 633 -3210 639 -2134
rect 593 -3222 639 -3210
rect -583 -3269 -341 -3263
rect -583 -3303 -571 -3269
rect -353 -3303 -341 -3269
rect -583 -3309 -341 -3303
rect -275 -3269 -33 -3263
rect -275 -3303 -263 -3269
rect -45 -3303 -33 -3269
rect -275 -3309 -33 -3303
rect 33 -3269 275 -3263
rect 33 -3303 45 -3269
rect 263 -3303 275 -3269
rect 33 -3309 275 -3303
rect 341 -3269 583 -3263
rect 341 -3303 353 -3269
rect 571 -3303 583 -3269
rect 341 -3309 583 -3303
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 5.5 l 1.25 m 5 nf 4 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 class mosfet compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1771420802
<< error_p >>
rect -918 3424 918 3436
rect -918 -3424 -906 3424
rect -882 3388 882 3400
rect -882 3284 -870 3388
rect -681 3328 -381 3331
rect -327 3328 -27 3331
rect 27 3328 327 3331
rect 381 3328 681 3331
rect -869 3284 -853 3300
rect -839 3284 -823 3300
rect -643 3293 -627 3309
rect -435 3293 -419 3309
rect -289 3293 -273 3309
rect -81 3293 -65 3309
rect 65 3293 81 3309
rect 273 3293 289 3309
rect 419 3293 435 3309
rect 627 3293 643 3309
rect -885 3268 -869 3284
rect -823 3268 -807 3284
rect -659 3277 -643 3293
rect -419 3277 -403 3293
rect -305 3277 -289 3293
rect -65 3277 -49 3293
rect 49 3277 65 3293
rect 289 3277 305 3293
rect 403 3277 419 3293
rect 643 3277 659 3293
rect 823 3284 839 3300
rect 853 3284 869 3300
rect 870 3284 882 3388
rect 807 3268 823 3284
rect 869 3268 885 3284
rect -882 -3268 -870 3268
rect -659 3261 -643 3263
rect -419 3261 -403 3263
rect -659 3247 -403 3261
rect -305 3261 -289 3263
rect -65 3261 -49 3263
rect -305 3247 -49 3261
rect 49 3261 65 3263
rect 289 3261 305 3263
rect 49 3247 305 3261
rect 403 3261 419 3263
rect 643 3261 659 3263
rect 403 3247 659 3261
rect -643 3231 -627 3247
rect -435 3231 -419 3247
rect -289 3231 -273 3247
rect -81 3231 -65 3247
rect 65 3231 81 3247
rect 273 3231 289 3247
rect 419 3231 435 3247
rect 627 3231 643 3247
rect -731 3201 -715 3217
rect -701 3201 -685 3217
rect -377 3201 -361 3217
rect -347 3201 -331 3217
rect -23 3201 -7 3217
rect 7 3201 23 3217
rect 331 3201 347 3217
rect 361 3201 377 3217
rect 685 3201 701 3217
rect 715 3201 731 3217
rect -747 3185 -731 3201
rect -685 3185 -669 3201
rect -393 3185 -377 3201
rect -331 3185 -315 3201
rect -39 3185 -23 3201
rect 23 3185 39 3201
rect 315 3185 331 3201
rect 377 3185 393 3201
rect 669 3185 685 3201
rect 731 3185 747 3201
rect -747 2127 -731 2143
rect -685 2127 -669 2143
rect -656 2127 -406 2128
rect -393 2127 -377 2143
rect -331 2127 -315 2143
rect -302 2127 -52 2128
rect -39 2127 -23 2143
rect 23 2127 39 2143
rect 52 2127 302 2128
rect 315 2127 331 2143
rect 377 2127 393 2143
rect 406 2127 656 2128
rect 669 2127 685 2143
rect 731 2127 747 2143
rect -731 2111 -715 2127
rect -701 2114 -361 2127
rect -701 2111 -685 2114
rect -377 2111 -361 2114
rect -347 2114 -7 2127
rect -347 2111 -331 2114
rect -23 2111 -7 2114
rect 7 2114 347 2127
rect 7 2111 23 2114
rect 331 2111 347 2114
rect 361 2114 701 2127
rect 361 2111 377 2114
rect 685 2111 701 2114
rect 715 2111 731 2127
rect -643 2081 -627 2097
rect -435 2081 -419 2097
rect -289 2081 -273 2097
rect -81 2081 -65 2097
rect 65 2081 81 2097
rect 273 2081 289 2097
rect 419 2081 435 2097
rect 627 2081 643 2097
rect -659 2065 -643 2081
rect -419 2065 -403 2081
rect -305 2065 -289 2081
rect -65 2065 -49 2081
rect 49 2065 65 2081
rect 289 2065 305 2081
rect 403 2065 419 2081
rect 643 2065 659 2081
rect -659 2035 -643 2051
rect -419 2035 -403 2051
rect -305 2035 -289 2051
rect -65 2035 -49 2051
rect 49 2035 65 2051
rect 289 2035 305 2051
rect 403 2035 419 2051
rect 643 2035 659 2051
rect -643 2019 -627 2035
rect -435 2019 -419 2035
rect -289 2019 -273 2035
rect -81 2019 -65 2035
rect 65 2019 81 2035
rect 273 2019 289 2035
rect 419 2019 435 2035
rect 627 2019 643 2035
rect -643 1961 -627 1977
rect -435 1961 -419 1977
rect -289 1961 -273 1977
rect -81 1961 -65 1977
rect 65 1961 81 1977
rect 273 1961 289 1977
rect 419 1961 435 1977
rect 627 1961 643 1977
rect -659 1945 -643 1961
rect -419 1945 -403 1961
rect -305 1945 -289 1961
rect -65 1945 -49 1961
rect 49 1945 65 1961
rect 289 1945 305 1961
rect 403 1945 419 1961
rect 643 1945 659 1961
rect -659 1929 -643 1931
rect -419 1929 -403 1931
rect -659 1915 -403 1929
rect -305 1929 -289 1931
rect -65 1929 -49 1931
rect -305 1915 -49 1929
rect 49 1929 65 1931
rect 289 1929 305 1931
rect 49 1915 305 1929
rect 403 1929 419 1931
rect 643 1929 659 1931
rect 403 1915 659 1929
rect -643 1899 -627 1915
rect -435 1899 -419 1915
rect -289 1899 -273 1915
rect -81 1899 -65 1915
rect 65 1899 81 1915
rect 273 1899 289 1915
rect 419 1899 435 1915
rect 627 1899 643 1915
rect -731 1869 -715 1885
rect -701 1869 -685 1885
rect -377 1869 -361 1885
rect -347 1869 -331 1885
rect -23 1869 -7 1885
rect 7 1869 23 1885
rect 331 1869 347 1885
rect 361 1869 377 1885
rect 685 1869 701 1885
rect 715 1869 731 1885
rect -747 1853 -731 1869
rect -685 1853 -669 1869
rect -393 1853 -377 1869
rect -331 1853 -315 1869
rect -39 1853 -23 1869
rect 23 1853 39 1869
rect 315 1853 331 1869
rect 377 1853 393 1869
rect 669 1853 685 1869
rect 731 1853 747 1869
rect -747 795 -731 811
rect -685 795 -669 811
rect -656 795 -406 796
rect -393 795 -377 811
rect -331 795 -315 811
rect -302 795 -52 796
rect -39 795 -23 811
rect 23 795 39 811
rect 52 795 302 796
rect 315 795 331 811
rect 377 795 393 811
rect 406 795 656 796
rect 669 795 685 811
rect 731 795 747 811
rect -731 779 -715 795
rect -701 782 -361 795
rect -701 779 -685 782
rect -377 779 -361 782
rect -347 782 -7 795
rect -347 779 -331 782
rect -23 779 -7 782
rect 7 782 347 795
rect 7 779 23 782
rect 331 779 347 782
rect 361 782 701 795
rect 361 779 377 782
rect 685 779 701 782
rect 715 779 731 795
rect -643 749 -627 765
rect -435 749 -419 765
rect -289 749 -273 765
rect -81 749 -65 765
rect 65 749 81 765
rect 273 749 289 765
rect 419 749 435 765
rect 627 749 643 765
rect -659 733 -643 749
rect -419 733 -403 749
rect -305 733 -289 749
rect -65 733 -49 749
rect 49 733 65 749
rect 289 733 305 749
rect 403 733 419 749
rect 643 733 659 749
rect -659 703 -643 719
rect -419 703 -403 719
rect -305 703 -289 719
rect -65 703 -49 719
rect 49 703 65 719
rect 289 703 305 719
rect 403 703 419 719
rect 643 703 659 719
rect -643 687 -627 703
rect -435 687 -419 703
rect -289 687 -273 703
rect -81 687 -65 703
rect 65 687 81 703
rect 273 687 289 703
rect 419 687 435 703
rect 627 687 643 703
rect -643 629 -627 645
rect -435 629 -419 645
rect -289 629 -273 645
rect -81 629 -65 645
rect 65 629 81 645
rect 273 629 289 645
rect 419 629 435 645
rect 627 629 643 645
rect -659 613 -643 629
rect -419 613 -403 629
rect -305 613 -289 629
rect -65 613 -49 629
rect 49 613 65 629
rect 289 613 305 629
rect 403 613 419 629
rect 643 613 659 629
rect -659 597 -643 599
rect -419 597 -403 599
rect -659 583 -403 597
rect -305 597 -289 599
rect -65 597 -49 599
rect -305 583 -49 597
rect 49 597 65 599
rect 289 597 305 599
rect 49 583 305 597
rect 403 597 419 599
rect 643 597 659 599
rect 403 583 659 597
rect -643 567 -627 583
rect -435 567 -419 583
rect -289 567 -273 583
rect -81 567 -65 583
rect 65 567 81 583
rect 273 567 289 583
rect 419 567 435 583
rect 627 567 643 583
rect -731 537 -715 553
rect -701 537 -685 553
rect -377 537 -361 553
rect -347 537 -331 553
rect -23 537 -7 553
rect 7 537 23 553
rect 331 537 347 553
rect 361 537 377 553
rect 685 537 701 553
rect 715 537 731 553
rect -747 521 -731 537
rect -685 521 -669 537
rect -393 521 -377 537
rect -331 521 -315 537
rect -39 521 -23 537
rect 23 521 39 537
rect 315 521 331 537
rect 377 521 393 537
rect 669 521 685 537
rect 731 521 747 537
rect -747 -537 -731 -521
rect -685 -537 -669 -521
rect -656 -537 -406 -536
rect -393 -537 -377 -521
rect -331 -537 -315 -521
rect -302 -537 -52 -536
rect -39 -537 -23 -521
rect 23 -537 39 -521
rect 52 -537 302 -536
rect 315 -537 331 -521
rect 377 -537 393 -521
rect 406 -537 656 -536
rect 669 -537 685 -521
rect 731 -537 747 -521
rect -731 -553 -715 -537
rect -701 -550 -361 -537
rect -701 -553 -685 -550
rect -377 -553 -361 -550
rect -347 -550 -7 -537
rect -347 -553 -331 -550
rect -23 -553 -7 -550
rect 7 -550 347 -537
rect 7 -553 23 -550
rect 331 -553 347 -550
rect 361 -550 701 -537
rect 361 -553 377 -550
rect 685 -553 701 -550
rect 715 -553 731 -537
rect -643 -583 -627 -567
rect -435 -583 -419 -567
rect -289 -583 -273 -567
rect -81 -583 -65 -567
rect 65 -583 81 -567
rect 273 -583 289 -567
rect 419 -583 435 -567
rect 627 -583 643 -567
rect -659 -599 -643 -583
rect -419 -599 -403 -583
rect -305 -599 -289 -583
rect -65 -599 -49 -583
rect 49 -599 65 -583
rect 289 -599 305 -583
rect 403 -599 419 -583
rect 643 -599 659 -583
rect -659 -629 -643 -613
rect -419 -629 -403 -613
rect -305 -629 -289 -613
rect -65 -629 -49 -613
rect 49 -629 65 -613
rect 289 -629 305 -613
rect 403 -629 419 -613
rect 643 -629 659 -613
rect -643 -645 -627 -629
rect -435 -645 -419 -629
rect -289 -645 -273 -629
rect -81 -645 -65 -629
rect 65 -645 81 -629
rect 273 -645 289 -629
rect 419 -645 435 -629
rect 627 -645 643 -629
rect -643 -703 -627 -687
rect -435 -703 -419 -687
rect -289 -703 -273 -687
rect -81 -703 -65 -687
rect 65 -703 81 -687
rect 273 -703 289 -687
rect 419 -703 435 -687
rect 627 -703 643 -687
rect -659 -719 -643 -703
rect -419 -719 -403 -703
rect -305 -719 -289 -703
rect -65 -719 -49 -703
rect 49 -719 65 -703
rect 289 -719 305 -703
rect 403 -719 419 -703
rect 643 -719 659 -703
rect -659 -735 -643 -733
rect -419 -735 -403 -733
rect -659 -749 -403 -735
rect -305 -735 -289 -733
rect -65 -735 -49 -733
rect -305 -749 -49 -735
rect 49 -735 65 -733
rect 289 -735 305 -733
rect 49 -749 305 -735
rect 403 -735 419 -733
rect 643 -735 659 -733
rect 403 -749 659 -735
rect -643 -765 -627 -749
rect -435 -765 -419 -749
rect -289 -765 -273 -749
rect -81 -765 -65 -749
rect 65 -765 81 -749
rect 273 -765 289 -749
rect 419 -765 435 -749
rect 627 -765 643 -749
rect -731 -795 -715 -779
rect -701 -795 -685 -779
rect -377 -795 -361 -779
rect -347 -795 -331 -779
rect -23 -795 -7 -779
rect 7 -795 23 -779
rect 331 -795 347 -779
rect 361 -795 377 -779
rect 685 -795 701 -779
rect 715 -795 731 -779
rect -747 -811 -731 -795
rect -685 -811 -669 -795
rect -393 -811 -377 -795
rect -331 -811 -315 -795
rect -39 -811 -23 -795
rect 23 -811 39 -795
rect 315 -811 331 -795
rect 377 -811 393 -795
rect 669 -811 685 -795
rect 731 -811 747 -795
rect -747 -1869 -731 -1853
rect -685 -1869 -669 -1853
rect -656 -1869 -406 -1868
rect -393 -1869 -377 -1853
rect -331 -1869 -315 -1853
rect -302 -1869 -52 -1868
rect -39 -1869 -23 -1853
rect 23 -1869 39 -1853
rect 52 -1869 302 -1868
rect 315 -1869 331 -1853
rect 377 -1869 393 -1853
rect 406 -1869 656 -1868
rect 669 -1869 685 -1853
rect 731 -1869 747 -1853
rect -731 -1885 -715 -1869
rect -701 -1882 -361 -1869
rect -701 -1885 -685 -1882
rect -377 -1885 -361 -1882
rect -347 -1882 -7 -1869
rect -347 -1885 -331 -1882
rect -23 -1885 -7 -1882
rect 7 -1882 347 -1869
rect 7 -1885 23 -1882
rect 331 -1885 347 -1882
rect 361 -1882 701 -1869
rect 361 -1885 377 -1882
rect 685 -1885 701 -1882
rect 715 -1885 731 -1869
rect -643 -1915 -627 -1899
rect -435 -1915 -419 -1899
rect -289 -1915 -273 -1899
rect -81 -1915 -65 -1899
rect 65 -1915 81 -1899
rect 273 -1915 289 -1899
rect 419 -1915 435 -1899
rect 627 -1915 643 -1899
rect -659 -1931 -643 -1915
rect -419 -1931 -403 -1915
rect -305 -1931 -289 -1915
rect -65 -1931 -49 -1915
rect 49 -1931 65 -1915
rect 289 -1931 305 -1915
rect 403 -1931 419 -1915
rect 643 -1931 659 -1915
rect -659 -1961 -643 -1945
rect -419 -1961 -403 -1945
rect -305 -1961 -289 -1945
rect -65 -1961 -49 -1945
rect 49 -1961 65 -1945
rect 289 -1961 305 -1945
rect 403 -1961 419 -1945
rect 643 -1961 659 -1945
rect -643 -1977 -627 -1961
rect -435 -1977 -419 -1961
rect -289 -1977 -273 -1961
rect -81 -1977 -65 -1961
rect 65 -1977 81 -1961
rect 273 -1977 289 -1961
rect 419 -1977 435 -1961
rect 627 -1977 643 -1961
rect -643 -2035 -627 -2019
rect -435 -2035 -419 -2019
rect -289 -2035 -273 -2019
rect -81 -2035 -65 -2019
rect 65 -2035 81 -2019
rect 273 -2035 289 -2019
rect 419 -2035 435 -2019
rect 627 -2035 643 -2019
rect -659 -2051 -643 -2035
rect -419 -2051 -403 -2035
rect -305 -2051 -289 -2035
rect -65 -2051 -49 -2035
rect 49 -2051 65 -2035
rect 289 -2051 305 -2035
rect 403 -2051 419 -2035
rect 643 -2051 659 -2035
rect -659 -2067 -643 -2065
rect -419 -2067 -403 -2065
rect -659 -2081 -403 -2067
rect -305 -2067 -289 -2065
rect -65 -2067 -49 -2065
rect -305 -2081 -49 -2067
rect 49 -2067 65 -2065
rect 289 -2067 305 -2065
rect 49 -2081 305 -2067
rect 403 -2067 419 -2065
rect 643 -2067 659 -2065
rect 403 -2081 659 -2067
rect -643 -2097 -627 -2081
rect -435 -2097 -419 -2081
rect -289 -2097 -273 -2081
rect -81 -2097 -65 -2081
rect 65 -2097 81 -2081
rect 273 -2097 289 -2081
rect 419 -2097 435 -2081
rect 627 -2097 643 -2081
rect -731 -2127 -715 -2111
rect -701 -2127 -685 -2111
rect -377 -2127 -361 -2111
rect -347 -2127 -331 -2111
rect -23 -2127 -7 -2111
rect 7 -2127 23 -2111
rect 331 -2127 347 -2111
rect 361 -2127 377 -2111
rect 685 -2127 701 -2111
rect 715 -2127 731 -2111
rect -747 -2143 -731 -2127
rect -685 -2143 -669 -2127
rect -393 -2143 -377 -2127
rect -331 -2143 -315 -2127
rect -39 -2143 -23 -2127
rect 23 -2143 39 -2127
rect 315 -2143 331 -2127
rect 377 -2143 393 -2127
rect 669 -2143 685 -2127
rect 731 -2143 747 -2127
rect -747 -3201 -731 -3185
rect -685 -3201 -669 -3185
rect -656 -3201 -406 -3200
rect -393 -3201 -377 -3185
rect -331 -3201 -315 -3185
rect -302 -3201 -52 -3200
rect -39 -3201 -23 -3185
rect 23 -3201 39 -3185
rect 52 -3201 302 -3200
rect 315 -3201 331 -3185
rect 377 -3201 393 -3185
rect 406 -3201 656 -3200
rect 669 -3201 685 -3185
rect 731 -3201 747 -3185
rect -731 -3217 -715 -3201
rect -701 -3214 -361 -3201
rect -701 -3217 -685 -3214
rect -377 -3217 -361 -3214
rect -347 -3214 -7 -3201
rect -347 -3217 -331 -3214
rect -23 -3217 -7 -3214
rect 7 -3214 347 -3201
rect 7 -3217 23 -3214
rect 331 -3217 347 -3214
rect 361 -3214 701 -3201
rect 361 -3217 377 -3214
rect 685 -3217 701 -3214
rect 715 -3217 731 -3201
rect -643 -3247 -627 -3231
rect -435 -3247 -419 -3231
rect -289 -3247 -273 -3231
rect -81 -3247 -65 -3231
rect 65 -3247 81 -3231
rect 273 -3247 289 -3231
rect 419 -3247 435 -3231
rect 627 -3247 643 -3231
rect -659 -3263 -643 -3247
rect -419 -3263 -403 -3247
rect -305 -3263 -289 -3247
rect -65 -3263 -49 -3247
rect 49 -3263 65 -3247
rect 289 -3263 305 -3247
rect 403 -3263 419 -3247
rect 643 -3263 659 -3247
rect 870 -3268 882 3268
rect -885 -3284 -869 -3268
rect -823 -3284 -807 -3268
rect -882 -3388 -870 -3284
rect -869 -3300 -853 -3284
rect -839 -3300 -823 -3284
rect -659 -3290 -643 -3277
rect -419 -3290 -403 -3277
rect -659 -3293 -403 -3290
rect -305 -3290 -289 -3277
rect -65 -3290 -49 -3277
rect -305 -3293 -49 -3290
rect 49 -3290 65 -3277
rect 289 -3290 305 -3277
rect 49 -3293 305 -3290
rect 403 -3290 419 -3277
rect 643 -3290 659 -3277
rect 807 -3284 823 -3268
rect 869 -3284 885 -3268
rect 403 -3293 659 -3290
rect -643 -3309 -627 -3293
rect -435 -3309 -419 -3293
rect -289 -3309 -273 -3293
rect -81 -3309 -65 -3293
rect 65 -3309 81 -3293
rect 273 -3309 289 -3293
rect 419 -3309 435 -3293
rect 627 -3309 643 -3293
rect 823 -3300 839 -3284
rect 853 -3300 869 -3284
rect 870 -3388 882 -3284
rect -882 -3400 882 -3388
rect 906 -3424 918 3424
rect -918 -3436 918 -3424
<< nwell >>
rect -906 -3424 906 3424
<< pmos >>
rect -656 2114 -406 3214
rect -302 2114 -52 3214
rect 52 2114 302 3214
rect 406 2114 656 3214
rect -656 782 -406 1882
rect -302 782 -52 1882
rect 52 782 302 1882
rect 406 782 656 1882
rect -656 -550 -406 550
rect -302 -550 -52 550
rect 52 -550 302 550
rect 406 -550 656 550
rect -656 -1882 -406 -782
rect -302 -1882 -52 -782
rect 52 -1882 302 -782
rect 406 -1882 656 -782
rect -656 -3214 -406 -2114
rect -302 -3214 -52 -2114
rect 52 -3214 302 -2114
rect 406 -3214 656 -2114
<< pdiff >>
rect -744 3201 -656 3214
rect -744 2127 -731 3201
rect -685 2127 -656 3201
rect -744 2114 -656 2127
rect -406 3201 -302 3214
rect -406 2127 -377 3201
rect -331 2127 -302 3201
rect -406 2114 -302 2127
rect -52 3201 52 3214
rect -52 2127 -23 3201
rect 23 2127 52 3201
rect -52 2114 52 2127
rect 302 3201 406 3214
rect 302 2127 331 3201
rect 377 2127 406 3201
rect 302 2114 406 2127
rect 656 3201 744 3214
rect 656 2127 685 3201
rect 731 2127 744 3201
rect 656 2114 744 2127
rect -744 1869 -656 1882
rect -744 795 -731 1869
rect -685 795 -656 1869
rect -744 782 -656 795
rect -406 1869 -302 1882
rect -406 795 -377 1869
rect -331 795 -302 1869
rect -406 782 -302 795
rect -52 1869 52 1882
rect -52 795 -23 1869
rect 23 795 52 1869
rect -52 782 52 795
rect 302 1869 406 1882
rect 302 795 331 1869
rect 377 795 406 1869
rect 302 782 406 795
rect 656 1869 744 1882
rect 656 795 685 1869
rect 731 795 744 1869
rect 656 782 744 795
rect -744 537 -656 550
rect -744 -537 -731 537
rect -685 -537 -656 537
rect -744 -550 -656 -537
rect -406 537 -302 550
rect -406 -537 -377 537
rect -331 -537 -302 537
rect -406 -550 -302 -537
rect -52 537 52 550
rect -52 -537 -23 537
rect 23 -537 52 537
rect -52 -550 52 -537
rect 302 537 406 550
rect 302 -537 331 537
rect 377 -537 406 537
rect 302 -550 406 -537
rect 656 537 744 550
rect 656 -537 685 537
rect 731 -537 744 537
rect 656 -550 744 -537
rect -744 -795 -656 -782
rect -744 -1869 -731 -795
rect -685 -1869 -656 -795
rect -744 -1882 -656 -1869
rect -406 -795 -302 -782
rect -406 -1869 -377 -795
rect -331 -1869 -302 -795
rect -406 -1882 -302 -1869
rect -52 -795 52 -782
rect -52 -1869 -23 -795
rect 23 -1869 52 -795
rect -52 -1882 52 -1869
rect 302 -795 406 -782
rect 302 -1869 331 -795
rect 377 -1869 406 -795
rect 302 -1882 406 -1869
rect 656 -795 744 -782
rect 656 -1869 685 -795
rect 731 -1869 744 -795
rect 656 -1882 744 -1869
rect -744 -2127 -656 -2114
rect -744 -3201 -731 -2127
rect -685 -3201 -656 -2127
rect -744 -3214 -656 -3201
rect -406 -2127 -302 -2114
rect -406 -3201 -377 -2127
rect -331 -3201 -302 -2127
rect -406 -3214 -302 -3201
rect -52 -2127 52 -2114
rect -52 -3201 -23 -2127
rect 23 -3201 52 -2127
rect -52 -3214 52 -3201
rect 302 -2127 406 -2114
rect 302 -3201 331 -2127
rect 377 -3201 406 -2127
rect 302 -3214 406 -3201
rect 656 -2127 744 -2114
rect 656 -3201 685 -2127
rect 731 -3201 744 -2127
rect 656 -3214 744 -3201
<< pdiffc >>
rect -731 2127 -685 3201
rect -377 2127 -331 3201
rect -23 2127 23 3201
rect 331 2127 377 3201
rect 685 2127 731 3201
rect -731 795 -685 1869
rect -377 795 -331 1869
rect -23 795 23 1869
rect 331 795 377 1869
rect 685 795 731 1869
rect -731 -537 -685 537
rect -377 -537 -331 537
rect -23 -537 23 537
rect 331 -537 377 537
rect 685 -537 731 537
rect -731 -1869 -685 -795
rect -377 -1869 -331 -795
rect -23 -1869 23 -795
rect 331 -1869 377 -795
rect 685 -1869 731 -795
rect -731 -3201 -685 -2127
rect -377 -3201 -331 -2127
rect -23 -3201 23 -2127
rect 331 -3201 377 -2127
rect 685 -3201 731 -2127
<< nsubdiff >>
rect -882 3328 882 3400
rect -882 3284 -810 3328
rect -882 -3284 -869 3284
rect -823 -3284 -810 3284
rect 810 3284 882 3328
rect -882 -3328 -810 -3284
rect 810 -3284 823 3284
rect 869 -3284 882 3284
rect 810 -3328 882 -3284
rect -882 -3400 882 -3328
<< nsubdiffcont >>
rect -869 -3284 -823 3284
rect 823 -3284 869 3284
<< poly >>
rect -656 3293 -406 3306
rect -656 3247 -643 3293
rect -419 3247 -406 3293
rect -656 3214 -406 3247
rect -302 3293 -52 3306
rect -302 3247 -289 3293
rect -65 3247 -52 3293
rect -302 3214 -52 3247
rect 52 3293 302 3306
rect 52 3247 65 3293
rect 289 3247 302 3293
rect 52 3214 302 3247
rect 406 3293 656 3306
rect 406 3247 419 3293
rect 643 3247 656 3293
rect 406 3214 656 3247
rect -656 2081 -406 2114
rect -656 2035 -643 2081
rect -419 2035 -406 2081
rect -656 2022 -406 2035
rect -302 2081 -52 2114
rect -302 2035 -289 2081
rect -65 2035 -52 2081
rect -302 2022 -52 2035
rect 52 2081 302 2114
rect 52 2035 65 2081
rect 289 2035 302 2081
rect 52 2022 302 2035
rect 406 2081 656 2114
rect 406 2035 419 2081
rect 643 2035 656 2081
rect 406 2022 656 2035
rect -656 1961 -406 1974
rect -656 1915 -643 1961
rect -419 1915 -406 1961
rect -656 1882 -406 1915
rect -302 1961 -52 1974
rect -302 1915 -289 1961
rect -65 1915 -52 1961
rect -302 1882 -52 1915
rect 52 1961 302 1974
rect 52 1915 65 1961
rect 289 1915 302 1961
rect 52 1882 302 1915
rect 406 1961 656 1974
rect 406 1915 419 1961
rect 643 1915 656 1961
rect 406 1882 656 1915
rect -656 749 -406 782
rect -656 703 -643 749
rect -419 703 -406 749
rect -656 690 -406 703
rect -302 749 -52 782
rect -302 703 -289 749
rect -65 703 -52 749
rect -302 690 -52 703
rect 52 749 302 782
rect 52 703 65 749
rect 289 703 302 749
rect 52 690 302 703
rect 406 749 656 782
rect 406 703 419 749
rect 643 703 656 749
rect 406 690 656 703
rect -656 629 -406 642
rect -656 583 -643 629
rect -419 583 -406 629
rect -656 550 -406 583
rect -302 629 -52 642
rect -302 583 -289 629
rect -65 583 -52 629
rect -302 550 -52 583
rect 52 629 302 642
rect 52 583 65 629
rect 289 583 302 629
rect 52 550 302 583
rect 406 629 656 642
rect 406 583 419 629
rect 643 583 656 629
rect 406 550 656 583
rect -656 -583 -406 -550
rect -656 -629 -643 -583
rect -419 -629 -406 -583
rect -656 -642 -406 -629
rect -302 -583 -52 -550
rect -302 -629 -289 -583
rect -65 -629 -52 -583
rect -302 -642 -52 -629
rect 52 -583 302 -550
rect 52 -629 65 -583
rect 289 -629 302 -583
rect 52 -642 302 -629
rect 406 -583 656 -550
rect 406 -629 419 -583
rect 643 -629 656 -583
rect 406 -642 656 -629
rect -656 -703 -406 -690
rect -656 -749 -643 -703
rect -419 -749 -406 -703
rect -656 -782 -406 -749
rect -302 -703 -52 -690
rect -302 -749 -289 -703
rect -65 -749 -52 -703
rect -302 -782 -52 -749
rect 52 -703 302 -690
rect 52 -749 65 -703
rect 289 -749 302 -703
rect 52 -782 302 -749
rect 406 -703 656 -690
rect 406 -749 419 -703
rect 643 -749 656 -703
rect 406 -782 656 -749
rect -656 -1915 -406 -1882
rect -656 -1961 -643 -1915
rect -419 -1961 -406 -1915
rect -656 -1974 -406 -1961
rect -302 -1915 -52 -1882
rect -302 -1961 -289 -1915
rect -65 -1961 -52 -1915
rect -302 -1974 -52 -1961
rect 52 -1915 302 -1882
rect 52 -1961 65 -1915
rect 289 -1961 302 -1915
rect 52 -1974 302 -1961
rect 406 -1915 656 -1882
rect 406 -1961 419 -1915
rect 643 -1961 656 -1915
rect 406 -1974 656 -1961
rect -656 -2035 -406 -2022
rect -656 -2081 -643 -2035
rect -419 -2081 -406 -2035
rect -656 -2114 -406 -2081
rect -302 -2035 -52 -2022
rect -302 -2081 -289 -2035
rect -65 -2081 -52 -2035
rect -302 -2114 -52 -2081
rect 52 -2035 302 -2022
rect 52 -2081 65 -2035
rect 289 -2081 302 -2035
rect 52 -2114 302 -2081
rect 406 -2035 656 -2022
rect 406 -2081 419 -2035
rect 643 -2081 656 -2035
rect 406 -2114 656 -2081
rect -656 -3247 -406 -3214
rect -656 -3293 -643 -3247
rect -419 -3293 -406 -3247
rect -656 -3306 -406 -3293
rect -302 -3247 -52 -3214
rect -302 -3293 -289 -3247
rect -65 -3293 -52 -3247
rect -302 -3306 -52 -3293
rect 52 -3247 302 -3214
rect 52 -3293 65 -3247
rect 289 -3293 302 -3247
rect 52 -3306 302 -3293
rect 406 -3247 656 -3214
rect 406 -3293 419 -3247
rect 643 -3293 656 -3247
rect 406 -3306 656 -3293
<< polycont >>
rect -643 3247 -419 3293
rect -289 3247 -65 3293
rect 65 3247 289 3293
rect 419 3247 643 3293
rect -643 2035 -419 2081
rect -289 2035 -65 2081
rect 65 2035 289 2081
rect 419 2035 643 2081
rect -643 1915 -419 1961
rect -289 1915 -65 1961
rect 65 1915 289 1961
rect 419 1915 643 1961
rect -643 703 -419 749
rect -289 703 -65 749
rect 65 703 289 749
rect 419 703 643 749
rect -643 583 -419 629
rect -289 583 -65 629
rect 65 583 289 629
rect 419 583 643 629
rect -643 -629 -419 -583
rect -289 -629 -65 -583
rect 65 -629 289 -583
rect 419 -629 643 -583
rect -643 -749 -419 -703
rect -289 -749 -65 -703
rect 65 -749 289 -703
rect 419 -749 643 -703
rect -643 -1961 -419 -1915
rect -289 -1961 -65 -1915
rect 65 -1961 289 -1915
rect 419 -1961 643 -1915
rect -643 -2081 -419 -2035
rect -289 -2081 -65 -2035
rect 65 -2081 289 -2035
rect 419 -2081 643 -2035
rect -643 -3293 -419 -3247
rect -289 -3293 -65 -3247
rect 65 -3293 289 -3247
rect 419 -3293 643 -3247
<< metal1 >>
rect -869 3341 869 3387
rect -869 -3341 -823 3341
rect -654 3247 -408 3293
rect -300 3247 -54 3293
rect 54 3247 300 3293
rect 408 3247 654 3293
rect -731 2116 -685 3212
rect -377 2116 -331 3212
rect -23 2116 23 3212
rect 331 2116 377 3212
rect 685 2116 731 3212
rect -654 2035 -408 2081
rect -300 2035 -54 2081
rect 54 2035 300 2081
rect 408 2035 654 2081
rect -654 1915 -408 1961
rect -300 1915 -54 1961
rect 54 1915 300 1961
rect 408 1915 654 1961
rect -731 784 -685 1880
rect -377 784 -331 1880
rect -23 784 23 1880
rect 331 784 377 1880
rect 685 784 731 1880
rect -654 703 -408 749
rect -300 703 -54 749
rect 54 703 300 749
rect 408 703 654 749
rect -654 583 -408 629
rect -300 583 -54 629
rect 54 583 300 629
rect 408 583 654 629
rect -731 -548 -685 548
rect -377 -548 -331 548
rect -23 -548 23 548
rect 331 -548 377 548
rect 685 -548 731 548
rect -654 -629 -408 -583
rect -300 -629 -54 -583
rect 54 -629 300 -583
rect 408 -629 654 -583
rect -654 -749 -408 -703
rect -300 -749 -54 -703
rect 54 -749 300 -703
rect 408 -749 654 -703
rect -731 -1880 -685 -784
rect -377 -1880 -331 -784
rect -23 -1880 23 -784
rect 331 -1880 377 -784
rect 685 -1880 731 -784
rect -654 -1961 -408 -1915
rect -300 -1961 -54 -1915
rect 54 -1961 300 -1915
rect 408 -1961 654 -1915
rect -654 -2081 -408 -2035
rect -300 -2081 -54 -2035
rect 54 -2081 300 -2035
rect 408 -2081 654 -2035
rect -731 -3212 -685 -2116
rect -377 -3212 -331 -2116
rect -23 -3212 23 -2116
rect 331 -3212 377 -2116
rect 685 -3212 731 -2116
rect -654 -3293 -408 -3247
rect -300 -3293 -54 -3247
rect 54 -3293 300 -3247
rect 408 -3293 654 -3247
rect 823 -3341 869 3341
rect -869 -3387 869 -3341
<< properties >>
string FIXED_BBOX -846 -3364 846 3364
string gencell pfet_03v3
string library gf180mcu
string parameters w 5.5 l 1.25 m 5 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 class mosfet full_metal 1 compatible {pfet_03v3 pfet_06v0}
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1771462974
<< error_p >>
rect -29 -132 29 -126
rect -29 -166 -17 -132
rect -29 -172 29 -166
<< nmos >>
rect -30 -94 30 156
<< ndiff >>
rect -88 144 -30 156
rect -88 -82 -76 144
rect -42 -82 -30 144
rect -88 -94 -30 -82
rect 30 144 88 156
rect 30 -82 42 144
rect 76 -82 88 144
rect 30 -94 88 -82
<< ndiffc >>
rect -76 -82 -42 144
rect 42 -82 76 144
<< poly >>
rect -30 156 30 182
rect -30 -116 30 -94
rect -33 -132 33 -116
rect -33 -166 -17 -132
rect 17 -166 33 -132
rect -33 -182 33 -166
<< polycont >>
rect -17 -166 17 -132
<< locali >>
rect -76 144 -42 160
rect -76 -98 -42 -82
rect 42 144 76 160
rect 42 -98 76 -82
rect -33 -166 -17 -132
rect 17 -166 33 -132
<< viali >>
rect -76 -82 -42 144
rect 42 -82 76 144
rect -17 -166 17 -132
<< metal1 >>
rect -82 144 -36 156
rect -82 -82 -76 144
rect -42 -82 -36 144
rect -82 -94 -36 -82
rect 36 144 82 156
rect 36 -82 42 144
rect 76 -82 82 144
rect 36 -94 82 -82
rect -29 -132 29 -126
rect -29 -166 -17 -132
rect 17 -166 29 -132
rect -29 -172 29 -166
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1.25 l 0.3 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 class mosfet compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

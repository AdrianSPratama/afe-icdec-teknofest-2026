magic
tech sky130A
magscale 1 2
timestamp 1771466212
<< nwell >>
rect -2440 140 5940 1440
rect 4060 -5440 5940 140
<< pwell >>
rect -2400 -3400 4000 100
<< psubdiff >>
rect -1500 80 -100 100
rect -1500 20 -1380 80
rect -220 20 -100 80
rect -1500 0 -100 20
rect -1500 -20 -1400 0
rect -2400 -120 -1600 -100
rect -2400 -180 -2280 -120
rect -1720 -180 -1600 -120
rect -2400 -200 -1600 -180
rect -2400 -220 -2300 -200
rect -2400 -780 -2380 -220
rect -2320 -780 -2300 -220
rect -2400 -800 -2300 -780
rect -1700 -220 -1600 -200
rect -1700 -780 -1680 -220
rect -1620 -780 -1600 -220
rect -1700 -800 -1600 -780
rect -2400 -820 -1600 -800
rect -2400 -880 -2280 -820
rect -1720 -880 -1600 -820
rect -2400 -900 -1600 -880
rect -1500 -1080 -1480 -20
rect -1420 -1080 -1400 -20
rect -1500 -1100 -1400 -1080
rect -200 -20 -100 0
rect -200 -1080 -180 -20
rect -120 -1080 -100 -20
rect -200 -1100 -100 -1080
rect -1500 -1120 -100 -1100
rect -1500 -1180 -1380 -1120
rect -220 -1180 -100 -1120
rect -1500 -1200 -100 -1180
rect 900 80 4000 100
rect 900 20 1020 80
rect 3880 20 4000 80
rect 900 0 4000 20
rect 900 -20 1000 0
rect -2400 -1320 -500 -1300
rect -2400 -1380 -2280 -1320
rect -620 -1380 -500 -1320
rect -2400 -1400 -500 -1380
rect -2400 -1420 -2300 -1400
rect -2400 -3280 -2380 -1420
rect -2320 -3280 -2300 -1420
rect -2400 -3300 -2300 -3280
rect -600 -1420 -500 -1400
rect -600 -3280 -580 -1420
rect -520 -3280 -500 -1420
rect 900 -1880 920 -20
rect 980 -1880 1000 -20
rect 3900 -20 4000 0
rect 1100 -120 1700 -100
rect 1100 -180 1160 -120
rect 1640 -180 1700 -120
rect 1100 -200 1700 -180
rect 1100 -800 1200 -200
rect 1600 -800 1700 -200
rect 1100 -900 1700 -800
rect 1800 -120 2400 -100
rect 1800 -180 1860 -120
rect 2340 -180 2400 -120
rect 1800 -200 2400 -180
rect 1800 -800 1900 -200
rect 2300 -800 2400 -200
rect 1800 -900 2400 -800
rect 2500 -120 3100 -100
rect 2500 -180 2560 -120
rect 3040 -180 3100 -120
rect 2500 -200 3100 -180
rect 2500 -800 2600 -200
rect 3000 -800 3100 -200
rect 2500 -900 3100 -800
rect 3200 -120 3800 -100
rect 3200 -180 3260 -120
rect 3740 -180 3800 -120
rect 3200 -200 3800 -180
rect 3200 -800 3300 -200
rect 3700 -800 3800 -200
rect 3200 -900 3800 -800
rect 1100 -1100 1700 -1000
rect 1100 -1700 1200 -1100
rect 1600 -1700 1700 -1100
rect 1100 -1720 1700 -1700
rect 1100 -1780 1160 -1720
rect 1640 -1780 1700 -1720
rect 1100 -1800 1700 -1780
rect 1800 -1100 2400 -1000
rect 1800 -1700 1900 -1100
rect 2300 -1700 2400 -1100
rect 1800 -1720 2400 -1700
rect 1800 -1780 1860 -1720
rect 2340 -1780 2400 -1720
rect 1800 -1800 2400 -1780
rect 2500 -1100 3100 -1000
rect 2500 -1700 2600 -1100
rect 3000 -1700 3100 -1100
rect 2500 -1720 3100 -1700
rect 2500 -1780 2560 -1720
rect 3040 -1780 3100 -1720
rect 2500 -1800 3100 -1780
rect 3200 -1100 3800 -1000
rect 3200 -1700 3300 -1100
rect 3700 -1700 3800 -1100
rect 3200 -1720 3800 -1700
rect 3200 -1780 3260 -1720
rect 3740 -1780 3800 -1720
rect 3200 -1800 3800 -1780
rect 900 -1900 1000 -1880
rect 3900 -1880 3920 -20
rect 3980 -1880 4000 -20
rect 3900 -1900 4000 -1880
rect 900 -1920 4000 -1900
rect 900 -1980 1020 -1920
rect 3880 -1980 4000 -1920
rect 900 -2000 4000 -1980
rect -600 -3300 -500 -3280
rect 900 -2120 1700 -2100
rect 900 -2180 1000 -2120
rect 1600 -2180 1700 -2120
rect 900 -2200 1700 -2180
rect 900 -2220 1000 -2200
rect 900 -3180 920 -2220
rect 980 -3180 1000 -2220
rect 900 -3200 1000 -3180
rect 1600 -2220 1700 -2200
rect 1600 -3180 1620 -2220
rect 1680 -3180 1700 -2220
rect 1600 -3200 1700 -3180
rect 900 -3220 1700 -3200
rect 900 -3280 1000 -3220
rect 1600 -3280 1700 -3220
rect 900 -3300 1700 -3280
rect 2300 -2120 4000 -2100
rect 2300 -2180 2420 -2120
rect 3880 -2180 4000 -2120
rect 2300 -2200 4000 -2180
rect 2300 -2220 2400 -2200
rect 2300 -3180 2320 -2220
rect 2380 -3180 2400 -2220
rect 2300 -3200 2400 -3180
rect 3900 -2220 4000 -2200
rect 3900 -3180 3920 -2220
rect 3980 -3180 4000 -2220
rect 3900 -3200 4000 -3180
rect 2300 -3220 4000 -3200
rect 2300 -3280 2420 -3220
rect 3880 -3280 4000 -3220
rect 2300 -3300 4000 -3280
rect -2400 -3320 -500 -3300
rect -2400 -3380 -2280 -3320
rect -620 -3380 -500 -3320
rect -2400 -3400 -500 -3380
<< nsubdiff >>
rect -2400 1380 800 1400
rect -2400 1320 -2280 1380
rect 680 1320 800 1380
rect -2400 1300 800 1320
rect -2400 1280 -2300 1300
rect -2400 320 -2380 1280
rect -2320 320 -2300 1280
rect -2400 300 -2300 320
rect 700 1280 800 1300
rect 700 320 720 1280
rect 780 320 800 1280
rect 700 300 800 320
rect -2400 280 800 300
rect -2400 220 -2280 280
rect 680 220 800 280
rect -2400 200 800 220
rect 900 1380 4000 1400
rect 900 1320 1020 1380
rect 3880 1320 4000 1380
rect 900 1300 4000 1320
rect 900 1280 1000 1300
rect 900 320 920 1280
rect 980 320 1000 1280
rect 900 300 1000 320
rect 3900 1280 4000 1300
rect 3900 320 3920 1280
rect 3980 320 4000 1280
rect 3900 300 4000 320
rect 900 280 4000 300
rect 900 220 1020 280
rect 3880 220 4000 280
rect 900 200 4000 220
rect 4100 1380 5900 1400
rect 4100 1320 4220 1380
rect 5780 1320 5900 1380
rect 4100 1300 5900 1320
rect 4100 1280 4200 1300
rect 4100 -5280 4120 1280
rect 4180 -5280 4200 1280
rect 4100 -5300 4200 -5280
rect 5800 1280 5900 1300
rect 5800 -5280 5820 1280
rect 5880 -5280 5900 1280
rect 5800 -5300 5900 -5280
rect 4100 -5320 5900 -5300
rect 4100 -5380 4220 -5320
rect 5780 -5380 5900 -5320
rect 4100 -5400 5900 -5380
<< psubdiffcont >>
rect -1380 20 -220 80
rect -2280 -180 -1720 -120
rect -2380 -780 -2320 -220
rect -1680 -780 -1620 -220
rect -2280 -880 -1720 -820
rect -1480 -1080 -1420 -20
rect -180 -1080 -120 -20
rect -1380 -1180 -220 -1120
rect 1020 20 3880 80
rect -2280 -1380 -620 -1320
rect -2380 -3280 -2320 -1420
rect -580 -3280 -520 -1420
rect 920 -1880 980 -20
rect 1160 -180 1640 -120
rect 1860 -180 2340 -120
rect 2560 -180 3040 -120
rect 3260 -180 3740 -120
rect 1160 -1780 1640 -1720
rect 1860 -1780 2340 -1720
rect 2560 -1780 3040 -1720
rect 3260 -1780 3740 -1720
rect 3920 -1880 3980 -20
rect 1020 -1980 3880 -1920
rect 1000 -2180 1600 -2120
rect 920 -3180 980 -2220
rect 1620 -3180 1680 -2220
rect 1000 -3280 1600 -3220
rect 2420 -2180 3880 -2120
rect 2320 -3180 2380 -2220
rect 3920 -3180 3980 -2220
rect 2420 -3280 3880 -3220
rect -2280 -3380 -620 -3320
<< nsubdiffcont >>
rect -2280 1320 680 1380
rect -2380 320 -2320 1280
rect 720 320 780 1280
rect -2280 220 680 280
rect 1020 1320 3880 1380
rect 920 320 980 1280
rect 3920 320 3980 1280
rect 1020 220 3880 280
rect 4220 1320 5780 1380
rect 4120 -5280 4180 1280
rect 5820 -5280 5880 1280
rect 4220 -5380 5780 -5320
<< locali >>
rect -2400 2080 -500 2100
rect -2400 2020 -2380 2080
rect -2320 2020 -2280 2080
rect -2220 2020 -2180 2080
rect -2120 2020 -2080 2080
rect -2020 2020 -1980 2080
rect -1920 2020 -1880 2080
rect -1820 2020 -1780 2080
rect -1720 2020 -1680 2080
rect -1620 2020 -1580 2080
rect -1520 2020 -1480 2080
rect -1420 2020 -1380 2080
rect -1320 2020 -1280 2080
rect -1220 2020 -1180 2080
rect -1120 2020 -1080 2080
rect -1020 2020 -980 2080
rect -920 2020 -880 2080
rect -820 2020 -780 2080
rect -720 2020 -680 2080
rect -620 2020 -580 2080
rect -520 2020 -500 2080
rect -2400 1980 -500 2020
rect -2400 1920 -2380 1980
rect -2320 1920 -2280 1980
rect -2220 1920 -2180 1980
rect -2120 1920 -2080 1980
rect -2020 1920 -1980 1980
rect -1920 1920 -1880 1980
rect -1820 1920 -1780 1980
rect -1720 1920 -1680 1980
rect -1620 1920 -1580 1980
rect -1520 1920 -1480 1980
rect -1420 1920 -1380 1980
rect -1320 1920 -1280 1980
rect -1220 1920 -1180 1980
rect -1120 1920 -1080 1980
rect -1020 1920 -980 1980
rect -920 1920 -880 1980
rect -820 1920 -780 1980
rect -720 1920 -680 1980
rect -620 1920 -580 1980
rect -520 1920 -500 1980
rect -2400 1880 -500 1920
rect -2400 1820 -2380 1880
rect -2320 1820 -2280 1880
rect -2220 1820 -2180 1880
rect -2120 1820 -2080 1880
rect -2020 1820 -1980 1880
rect -1920 1820 -1880 1880
rect -1820 1820 -1780 1880
rect -1720 1820 -1680 1880
rect -1620 1820 -1580 1880
rect -1520 1820 -1480 1880
rect -1420 1820 -1380 1880
rect -1320 1820 -1280 1880
rect -1220 1820 -1180 1880
rect -1120 1820 -1080 1880
rect -1020 1820 -980 1880
rect -920 1820 -880 1880
rect -820 1820 -780 1880
rect -720 1820 -680 1880
rect -620 1820 -580 1880
rect -520 1820 -500 1880
rect -2400 1780 -500 1820
rect -2400 1720 -2380 1780
rect -2320 1720 -2280 1780
rect -2220 1720 -2180 1780
rect -2120 1720 -2080 1780
rect -2020 1720 -1980 1780
rect -1920 1720 -1880 1780
rect -1820 1720 -1780 1780
rect -1720 1720 -1680 1780
rect -1620 1720 -1580 1780
rect -1520 1720 -1480 1780
rect -1420 1720 -1380 1780
rect -1320 1720 -1280 1780
rect -1220 1720 -1180 1780
rect -1120 1720 -1080 1780
rect -1020 1720 -980 1780
rect -920 1720 -880 1780
rect -820 1720 -780 1780
rect -720 1720 -680 1780
rect -620 1720 -580 1780
rect -520 1720 -500 1780
rect -2400 1680 -500 1720
rect -2400 1620 -2380 1680
rect -2320 1620 -2280 1680
rect -2220 1620 -2180 1680
rect -2120 1620 -2080 1680
rect -2020 1620 -1980 1680
rect -1920 1620 -1880 1680
rect -1820 1620 -1780 1680
rect -1720 1620 -1680 1680
rect -1620 1620 -1580 1680
rect -1520 1620 -1480 1680
rect -1420 1620 -1380 1680
rect -1320 1620 -1280 1680
rect -1220 1620 -1180 1680
rect -1120 1620 -1080 1680
rect -1020 1620 -980 1680
rect -920 1620 -880 1680
rect -820 1620 -780 1680
rect -720 1620 -680 1680
rect -620 1620 -580 1680
rect -520 1620 -500 1680
rect -2400 1580 -500 1620
rect -2400 1520 -2380 1580
rect -2320 1520 -2280 1580
rect -2220 1520 -2180 1580
rect -2120 1520 -2080 1580
rect -2020 1520 -1980 1580
rect -1920 1520 -1880 1580
rect -1820 1520 -1780 1580
rect -1720 1520 -1680 1580
rect -1620 1520 -1580 1580
rect -1520 1520 -1480 1580
rect -1420 1520 -1380 1580
rect -1320 1520 -1280 1580
rect -1220 1520 -1180 1580
rect -1120 1520 -1080 1580
rect -1020 1520 -980 1580
rect -920 1520 -880 1580
rect -820 1520 -780 1580
rect -720 1520 -680 1580
rect -620 1520 -580 1580
rect -520 1520 -500 1580
rect -2400 1480 -500 1520
rect -2400 1420 -2380 1480
rect -2320 1420 -2280 1480
rect -2220 1420 -2180 1480
rect -2120 1420 -2080 1480
rect -2020 1420 -1980 1480
rect -1920 1420 -1880 1480
rect -1820 1420 -1780 1480
rect -1720 1420 -1680 1480
rect -1620 1420 -1580 1480
rect -1520 1420 -1480 1480
rect -1420 1420 -1380 1480
rect -1320 1420 -1280 1480
rect -1220 1420 -1180 1480
rect -1120 1420 -1080 1480
rect -1020 1420 -980 1480
rect -920 1420 -880 1480
rect -820 1420 -780 1480
rect -720 1420 -680 1480
rect -620 1420 -580 1480
rect -520 1420 -500 1480
rect -2400 1400 -500 1420
rect -2400 1380 5900 1400
rect -2400 1320 -2280 1380
rect 680 1320 1020 1380
rect 3880 1320 4220 1380
rect 5780 1320 5900 1380
rect -2400 1300 5900 1320
rect -2400 1280 -2300 1300
rect -2400 320 -2380 1280
rect -2320 320 -2300 1280
rect -1880 520 -1780 1300
rect -1260 520 -1160 1300
rect -480 520 -380 1300
rect 140 520 240 1300
rect 700 1280 1000 1300
rect -2400 300 -2300 320
rect 700 320 720 1280
rect 780 320 920 1280
rect 980 320 1000 1280
rect 1500 600 1600 1300
rect 2100 600 2200 1300
rect 2700 600 2800 1300
rect 3300 600 3400 1300
rect 3900 1280 4200 1300
rect 700 300 1000 320
rect 3900 320 3920 1280
rect 3980 320 4120 1280
rect 3900 300 4120 320
rect -2400 280 4120 300
rect -2400 220 -2280 280
rect 680 220 1020 280
rect 3880 220 4120 280
rect -2400 200 4120 220
rect -2400 80 4000 100
rect -2400 20 -1380 80
rect -220 20 1020 80
rect 3880 20 4000 80
rect -2400 0 4000 20
rect -2400 -20 -1400 0
rect -2400 -120 -1480 -20
rect -2400 -180 -2280 -120
rect -1720 -180 -1480 -120
rect -2400 -200 -1480 -180
rect -2400 -220 -2300 -200
rect -2400 -780 -2380 -220
rect -2320 -780 -2300 -220
rect -2400 -800 -2300 -780
rect -1700 -220 -1480 -200
rect -1700 -780 -1680 -220
rect -1620 -780 -1480 -220
rect -1700 -800 -1480 -780
rect -2400 -820 -1480 -800
rect -2400 -880 -2280 -820
rect -1720 -880 -1480 -820
rect -2400 -1080 -1480 -880
rect -1420 -1080 -1400 -20
rect -980 -900 -880 0
rect -200 -20 4000 0
rect -2400 -1100 -1400 -1080
rect -200 -1080 -180 -20
rect -120 -1080 920 -20
rect -200 -1100 920 -1080
rect -2400 -1120 920 -1100
rect -2400 -1180 -1380 -1120
rect -220 -1180 920 -1120
rect -2400 -1320 920 -1180
rect -2400 -1380 -2280 -1320
rect -620 -1380 920 -1320
rect -2400 -1400 920 -1380
rect -2400 -1420 -2300 -1400
rect -2400 -3280 -2380 -1420
rect -2320 -3280 -2300 -1420
rect -2400 -3300 -2300 -3280
rect -600 -1420 920 -1400
rect -600 -3280 -580 -1420
rect -520 -1880 920 -1420
rect 980 -60 3920 -20
rect 980 -1840 1060 -60
rect 1140 -120 1660 -60
rect 1140 -180 1160 -120
rect 1640 -180 1660 -120
rect 1140 -200 1660 -180
rect 1700 -900 1800 -100
rect 1840 -120 2360 -60
rect 1840 -180 1860 -120
rect 2340 -180 2360 -120
rect 1840 -200 2360 -180
rect 2400 -120 2500 -100
rect 2400 -180 2420 -120
rect 2480 -180 2500 -120
rect 2400 -220 2500 -180
rect 2540 -120 3060 -60
rect 2540 -180 2560 -120
rect 3040 -180 3060 -120
rect 2540 -200 3060 -180
rect 2400 -280 2420 -220
rect 2480 -280 2500 -220
rect 2400 -320 2500 -280
rect 2400 -380 2420 -320
rect 2480 -380 2500 -320
rect 2400 -420 2500 -380
rect 2400 -480 2420 -420
rect 2480 -480 2500 -420
rect 2400 -520 2500 -480
rect 2400 -580 2420 -520
rect 2480 -580 2500 -520
rect 2400 -620 2500 -580
rect 2400 -680 2420 -620
rect 2480 -680 2500 -620
rect 2400 -900 2500 -680
rect 3100 -900 3200 -100
rect 3240 -120 3760 -60
rect 3240 -180 3260 -120
rect 3740 -180 3760 -120
rect 3240 -200 3760 -180
rect 1100 -1000 3800 -900
rect 1140 -1720 1660 -1700
rect 1140 -1780 1160 -1720
rect 1640 -1780 1660 -1720
rect 1140 -1840 1660 -1780
rect 1700 -1800 1800 -1000
rect 2400 -1220 2500 -1000
rect 2400 -1280 2420 -1220
rect 2480 -1280 2500 -1220
rect 2400 -1320 2500 -1280
rect 2400 -1380 2420 -1320
rect 2480 -1380 2500 -1320
rect 2400 -1420 2500 -1380
rect 2400 -1480 2420 -1420
rect 2480 -1480 2500 -1420
rect 2400 -1520 2500 -1480
rect 2400 -1580 2420 -1520
rect 2480 -1580 2500 -1520
rect 2400 -1620 2500 -1580
rect 2400 -1680 2420 -1620
rect 2480 -1680 2500 -1620
rect 1840 -1720 2360 -1700
rect 1840 -1780 1860 -1720
rect 2340 -1780 2360 -1720
rect 1840 -1840 2360 -1780
rect 2400 -1720 2500 -1680
rect 2400 -1780 2420 -1720
rect 2480 -1780 2500 -1720
rect 2400 -1800 2500 -1780
rect 2540 -1720 3060 -1700
rect 2540 -1780 2560 -1720
rect 3040 -1780 3060 -1720
rect 2540 -1840 3060 -1780
rect 3100 -1800 3200 -1000
rect 3240 -1720 3760 -1700
rect 3240 -1780 3260 -1720
rect 3740 -1780 3760 -1720
rect 3240 -1840 3760 -1780
rect 3840 -1840 3920 -60
rect 980 -1880 3920 -1840
rect 3980 -1880 4000 -20
rect -520 -1920 4000 -1880
rect -520 -1980 1020 -1920
rect 3880 -1980 4000 -1920
rect -520 -2120 4000 -1980
rect -520 -2180 1000 -2120
rect 1600 -2180 2420 -2120
rect 3880 -2180 4000 -2120
rect -520 -2200 4000 -2180
rect -520 -2220 1000 -2200
rect -520 -3180 920 -2220
rect 980 -3180 1000 -2220
rect 1600 -2220 2400 -2200
rect -520 -3200 1000 -3180
rect 1040 -3200 1140 -2400
rect 1600 -3180 1620 -2220
rect 1680 -3180 2320 -2220
rect 2380 -3180 2400 -2220
rect 3900 -2220 4000 -2200
rect 1600 -3200 2400 -3180
rect 2780 -3200 2880 -2500
rect 3400 -3200 3500 -2500
rect 3900 -3180 3920 -2220
rect 3980 -3180 4000 -2220
rect 3900 -3200 4000 -3180
rect -520 -3220 4000 -3200
rect -520 -3280 1000 -3220
rect 1600 -3280 2420 -3220
rect 3880 -3280 4000 -3220
rect -600 -3300 4000 -3280
rect -2400 -3320 4000 -3300
rect -2400 -3380 -2280 -3320
rect -620 -3380 4000 -3320
rect -2400 -3400 4000 -3380
rect -2400 -3420 -500 -3400
rect -2400 -3480 -2380 -3420
rect -2320 -3480 -2280 -3420
rect -2220 -3480 -2180 -3420
rect -2120 -3480 -2080 -3420
rect -2020 -3480 -1980 -3420
rect -1920 -3480 -1880 -3420
rect -1820 -3480 -1780 -3420
rect -1720 -3480 -1680 -3420
rect -1620 -3480 -1580 -3420
rect -1520 -3480 -1480 -3420
rect -1420 -3480 -1380 -3420
rect -1320 -3480 -1280 -3420
rect -1220 -3480 -1180 -3420
rect -1120 -3480 -1080 -3420
rect -1020 -3480 -980 -3420
rect -920 -3480 -880 -3420
rect -820 -3480 -780 -3420
rect -720 -3480 -680 -3420
rect -620 -3480 -580 -3420
rect -520 -3480 -500 -3420
rect -2400 -3520 -500 -3480
rect -2400 -3580 -2380 -3520
rect -2320 -3580 -2280 -3520
rect -2220 -3580 -2180 -3520
rect -2120 -3580 -2080 -3520
rect -2020 -3580 -1980 -3520
rect -1920 -3580 -1880 -3520
rect -1820 -3580 -1780 -3520
rect -1720 -3580 -1680 -3520
rect -1620 -3580 -1580 -3520
rect -1520 -3580 -1480 -3520
rect -1420 -3580 -1380 -3520
rect -1320 -3580 -1280 -3520
rect -1220 -3580 -1180 -3520
rect -1120 -3580 -1080 -3520
rect -1020 -3580 -980 -3520
rect -920 -3580 -880 -3520
rect -820 -3580 -780 -3520
rect -720 -3580 -680 -3520
rect -620 -3580 -580 -3520
rect -520 -3580 -500 -3520
rect -2400 -3620 -500 -3580
rect -2400 -3680 -2380 -3620
rect -2320 -3680 -2280 -3620
rect -2220 -3680 -2180 -3620
rect -2120 -3680 -2080 -3620
rect -2020 -3680 -1980 -3620
rect -1920 -3680 -1880 -3620
rect -1820 -3680 -1780 -3620
rect -1720 -3680 -1680 -3620
rect -1620 -3680 -1580 -3620
rect -1520 -3680 -1480 -3620
rect -1420 -3680 -1380 -3620
rect -1320 -3680 -1280 -3620
rect -1220 -3680 -1180 -3620
rect -1120 -3680 -1080 -3620
rect -1020 -3680 -980 -3620
rect -920 -3680 -880 -3620
rect -820 -3680 -780 -3620
rect -720 -3680 -680 -3620
rect -620 -3680 -580 -3620
rect -520 -3680 -500 -3620
rect -2400 -3720 -500 -3680
rect -2400 -3780 -2380 -3720
rect -2320 -3780 -2280 -3720
rect -2220 -3780 -2180 -3720
rect -2120 -3780 -2080 -3720
rect -2020 -3780 -1980 -3720
rect -1920 -3780 -1880 -3720
rect -1820 -3780 -1780 -3720
rect -1720 -3780 -1680 -3720
rect -1620 -3780 -1580 -3720
rect -1520 -3780 -1480 -3720
rect -1420 -3780 -1380 -3720
rect -1320 -3780 -1280 -3720
rect -1220 -3780 -1180 -3720
rect -1120 -3780 -1080 -3720
rect -1020 -3780 -980 -3720
rect -920 -3780 -880 -3720
rect -820 -3780 -780 -3720
rect -720 -3780 -680 -3720
rect -620 -3780 -580 -3720
rect -520 -3780 -500 -3720
rect -2400 -3820 -500 -3780
rect -2400 -3880 -2380 -3820
rect -2320 -3880 -2280 -3820
rect -2220 -3880 -2180 -3820
rect -2120 -3880 -2080 -3820
rect -2020 -3880 -1980 -3820
rect -1920 -3880 -1880 -3820
rect -1820 -3880 -1780 -3820
rect -1720 -3880 -1680 -3820
rect -1620 -3880 -1580 -3820
rect -1520 -3880 -1480 -3820
rect -1420 -3880 -1380 -3820
rect -1320 -3880 -1280 -3820
rect -1220 -3880 -1180 -3820
rect -1120 -3880 -1080 -3820
rect -1020 -3880 -980 -3820
rect -920 -3880 -880 -3820
rect -820 -3880 -780 -3820
rect -720 -3880 -680 -3820
rect -620 -3880 -580 -3820
rect -520 -3880 -500 -3820
rect -2400 -3920 -500 -3880
rect -2400 -3980 -2380 -3920
rect -2320 -3980 -2280 -3920
rect -2220 -3980 -2180 -3920
rect -2120 -3980 -2080 -3920
rect -2020 -3980 -1980 -3920
rect -1920 -3980 -1880 -3920
rect -1820 -3980 -1780 -3920
rect -1720 -3980 -1680 -3920
rect -1620 -3980 -1580 -3920
rect -1520 -3980 -1480 -3920
rect -1420 -3980 -1380 -3920
rect -1320 -3980 -1280 -3920
rect -1220 -3980 -1180 -3920
rect -1120 -3980 -1080 -3920
rect -1020 -3980 -980 -3920
rect -920 -3980 -880 -3920
rect -820 -3980 -780 -3920
rect -720 -3980 -680 -3920
rect -620 -3980 -580 -3920
rect -520 -3980 -500 -3920
rect -2400 -4020 -500 -3980
rect -2400 -4080 -2380 -4020
rect -2320 -4080 -2280 -4020
rect -2220 -4080 -2180 -4020
rect -2120 -4080 -2080 -4020
rect -2020 -4080 -1980 -4020
rect -1920 -4080 -1880 -4020
rect -1820 -4080 -1780 -4020
rect -1720 -4080 -1680 -4020
rect -1620 -4080 -1580 -4020
rect -1520 -4080 -1480 -4020
rect -1420 -4080 -1380 -4020
rect -1320 -4080 -1280 -4020
rect -1220 -4080 -1180 -4020
rect -1120 -4080 -1080 -4020
rect -1020 -4080 -980 -4020
rect -920 -4080 -880 -4020
rect -820 -4080 -780 -4020
rect -720 -4080 -680 -4020
rect -620 -4080 -580 -4020
rect -520 -4080 -500 -4020
rect -2400 -4100 -500 -4080
rect 4100 -5280 4120 200
rect 4180 -5280 4200 1280
rect 4100 -5300 4200 -5280
rect 4620 -5300 4720 1300
rect 5240 -5300 5340 1300
rect 5800 1280 5900 1300
rect 5800 -5280 5820 1280
rect 5880 -5280 5900 1280
rect 5800 -5300 5900 -5280
rect 4100 -5320 5900 -5300
rect 4100 -5380 4220 -5320
rect 5780 -5380 5900 -5320
rect 4100 -5400 5900 -5380
<< viali >>
rect -2380 2020 -2320 2080
rect -2280 2020 -2220 2080
rect -2180 2020 -2120 2080
rect -2080 2020 -2020 2080
rect -1980 2020 -1920 2080
rect -1880 2020 -1820 2080
rect -1780 2020 -1720 2080
rect -1680 2020 -1620 2080
rect -1580 2020 -1520 2080
rect -1480 2020 -1420 2080
rect -1380 2020 -1320 2080
rect -1280 2020 -1220 2080
rect -1180 2020 -1120 2080
rect -1080 2020 -1020 2080
rect -980 2020 -920 2080
rect -880 2020 -820 2080
rect -780 2020 -720 2080
rect -680 2020 -620 2080
rect -580 2020 -520 2080
rect -2380 1920 -2320 1980
rect -2280 1920 -2220 1980
rect -2180 1920 -2120 1980
rect -2080 1920 -2020 1980
rect -1980 1920 -1920 1980
rect -1880 1920 -1820 1980
rect -1780 1920 -1720 1980
rect -1680 1920 -1620 1980
rect -1580 1920 -1520 1980
rect -1480 1920 -1420 1980
rect -1380 1920 -1320 1980
rect -1280 1920 -1220 1980
rect -1180 1920 -1120 1980
rect -1080 1920 -1020 1980
rect -980 1920 -920 1980
rect -880 1920 -820 1980
rect -780 1920 -720 1980
rect -680 1920 -620 1980
rect -580 1920 -520 1980
rect -2380 1820 -2320 1880
rect -2280 1820 -2220 1880
rect -2180 1820 -2120 1880
rect -2080 1820 -2020 1880
rect -1980 1820 -1920 1880
rect -1880 1820 -1820 1880
rect -1780 1820 -1720 1880
rect -1680 1820 -1620 1880
rect -1580 1820 -1520 1880
rect -1480 1820 -1420 1880
rect -1380 1820 -1320 1880
rect -1280 1820 -1220 1880
rect -1180 1820 -1120 1880
rect -1080 1820 -1020 1880
rect -980 1820 -920 1880
rect -880 1820 -820 1880
rect -780 1820 -720 1880
rect -680 1820 -620 1880
rect -580 1820 -520 1880
rect -2380 1720 -2320 1780
rect -2280 1720 -2220 1780
rect -2180 1720 -2120 1780
rect -2080 1720 -2020 1780
rect -1980 1720 -1920 1780
rect -1880 1720 -1820 1780
rect -1780 1720 -1720 1780
rect -1680 1720 -1620 1780
rect -1580 1720 -1520 1780
rect -1480 1720 -1420 1780
rect -1380 1720 -1320 1780
rect -1280 1720 -1220 1780
rect -1180 1720 -1120 1780
rect -1080 1720 -1020 1780
rect -980 1720 -920 1780
rect -880 1720 -820 1780
rect -780 1720 -720 1780
rect -680 1720 -620 1780
rect -580 1720 -520 1780
rect -2380 1620 -2320 1680
rect -2280 1620 -2220 1680
rect -2180 1620 -2120 1680
rect -2080 1620 -2020 1680
rect -1980 1620 -1920 1680
rect -1880 1620 -1820 1680
rect -1780 1620 -1720 1680
rect -1680 1620 -1620 1680
rect -1580 1620 -1520 1680
rect -1480 1620 -1420 1680
rect -1380 1620 -1320 1680
rect -1280 1620 -1220 1680
rect -1180 1620 -1120 1680
rect -1080 1620 -1020 1680
rect -980 1620 -920 1680
rect -880 1620 -820 1680
rect -780 1620 -720 1680
rect -680 1620 -620 1680
rect -580 1620 -520 1680
rect -2380 1520 -2320 1580
rect -2280 1520 -2220 1580
rect -2180 1520 -2120 1580
rect -2080 1520 -2020 1580
rect -1980 1520 -1920 1580
rect -1880 1520 -1820 1580
rect -1780 1520 -1720 1580
rect -1680 1520 -1620 1580
rect -1580 1520 -1520 1580
rect -1480 1520 -1420 1580
rect -1380 1520 -1320 1580
rect -1280 1520 -1220 1580
rect -1180 1520 -1120 1580
rect -1080 1520 -1020 1580
rect -980 1520 -920 1580
rect -880 1520 -820 1580
rect -780 1520 -720 1580
rect -680 1520 -620 1580
rect -580 1520 -520 1580
rect -2380 1420 -2320 1480
rect -2280 1420 -2220 1480
rect -2180 1420 -2120 1480
rect -2080 1420 -2020 1480
rect -1980 1420 -1920 1480
rect -1880 1420 -1820 1480
rect -1780 1420 -1720 1480
rect -1680 1420 -1620 1480
rect -1580 1420 -1520 1480
rect -1480 1420 -1420 1480
rect -1380 1420 -1320 1480
rect -1280 1420 -1220 1480
rect -1180 1420 -1120 1480
rect -1080 1420 -1020 1480
rect -980 1420 -920 1480
rect -880 1420 -820 1480
rect -780 1420 -720 1480
rect -680 1420 -620 1480
rect -580 1420 -520 1480
rect 2420 -180 2480 -120
rect 2420 -280 2480 -220
rect 2420 -380 2480 -320
rect 2420 -480 2480 -420
rect 2420 -580 2480 -520
rect 2420 -680 2480 -620
rect 2420 -1280 2480 -1220
rect 2420 -1380 2480 -1320
rect 2420 -1480 2480 -1420
rect 2420 -1580 2480 -1520
rect 2420 -1680 2480 -1620
rect 2420 -1780 2480 -1720
rect -2380 -3480 -2320 -3420
rect -2280 -3480 -2220 -3420
rect -2180 -3480 -2120 -3420
rect -2080 -3480 -2020 -3420
rect -1980 -3480 -1920 -3420
rect -1880 -3480 -1820 -3420
rect -1780 -3480 -1720 -3420
rect -1680 -3480 -1620 -3420
rect -1580 -3480 -1520 -3420
rect -1480 -3480 -1420 -3420
rect -1380 -3480 -1320 -3420
rect -1280 -3480 -1220 -3420
rect -1180 -3480 -1120 -3420
rect -1080 -3480 -1020 -3420
rect -980 -3480 -920 -3420
rect -880 -3480 -820 -3420
rect -780 -3480 -720 -3420
rect -680 -3480 -620 -3420
rect -580 -3480 -520 -3420
rect -2380 -3580 -2320 -3520
rect -2280 -3580 -2220 -3520
rect -2180 -3580 -2120 -3520
rect -2080 -3580 -2020 -3520
rect -1980 -3580 -1920 -3520
rect -1880 -3580 -1820 -3520
rect -1780 -3580 -1720 -3520
rect -1680 -3580 -1620 -3520
rect -1580 -3580 -1520 -3520
rect -1480 -3580 -1420 -3520
rect -1380 -3580 -1320 -3520
rect -1280 -3580 -1220 -3520
rect -1180 -3580 -1120 -3520
rect -1080 -3580 -1020 -3520
rect -980 -3580 -920 -3520
rect -880 -3580 -820 -3520
rect -780 -3580 -720 -3520
rect -680 -3580 -620 -3520
rect -580 -3580 -520 -3520
rect -2380 -3680 -2320 -3620
rect -2280 -3680 -2220 -3620
rect -2180 -3680 -2120 -3620
rect -2080 -3680 -2020 -3620
rect -1980 -3680 -1920 -3620
rect -1880 -3680 -1820 -3620
rect -1780 -3680 -1720 -3620
rect -1680 -3680 -1620 -3620
rect -1580 -3680 -1520 -3620
rect -1480 -3680 -1420 -3620
rect -1380 -3680 -1320 -3620
rect -1280 -3680 -1220 -3620
rect -1180 -3680 -1120 -3620
rect -1080 -3680 -1020 -3620
rect -980 -3680 -920 -3620
rect -880 -3680 -820 -3620
rect -780 -3680 -720 -3620
rect -680 -3680 -620 -3620
rect -580 -3680 -520 -3620
rect -2380 -3780 -2320 -3720
rect -2280 -3780 -2220 -3720
rect -2180 -3780 -2120 -3720
rect -2080 -3780 -2020 -3720
rect -1980 -3780 -1920 -3720
rect -1880 -3780 -1820 -3720
rect -1780 -3780 -1720 -3720
rect -1680 -3780 -1620 -3720
rect -1580 -3780 -1520 -3720
rect -1480 -3780 -1420 -3720
rect -1380 -3780 -1320 -3720
rect -1280 -3780 -1220 -3720
rect -1180 -3780 -1120 -3720
rect -1080 -3780 -1020 -3720
rect -980 -3780 -920 -3720
rect -880 -3780 -820 -3720
rect -780 -3780 -720 -3720
rect -680 -3780 -620 -3720
rect -580 -3780 -520 -3720
rect -2380 -3880 -2320 -3820
rect -2280 -3880 -2220 -3820
rect -2180 -3880 -2120 -3820
rect -2080 -3880 -2020 -3820
rect -1980 -3880 -1920 -3820
rect -1880 -3880 -1820 -3820
rect -1780 -3880 -1720 -3820
rect -1680 -3880 -1620 -3820
rect -1580 -3880 -1520 -3820
rect -1480 -3880 -1420 -3820
rect -1380 -3880 -1320 -3820
rect -1280 -3880 -1220 -3820
rect -1180 -3880 -1120 -3820
rect -1080 -3880 -1020 -3820
rect -980 -3880 -920 -3820
rect -880 -3880 -820 -3820
rect -780 -3880 -720 -3820
rect -680 -3880 -620 -3820
rect -580 -3880 -520 -3820
rect -2380 -3980 -2320 -3920
rect -2280 -3980 -2220 -3920
rect -2180 -3980 -2120 -3920
rect -2080 -3980 -2020 -3920
rect -1980 -3980 -1920 -3920
rect -1880 -3980 -1820 -3920
rect -1780 -3980 -1720 -3920
rect -1680 -3980 -1620 -3920
rect -1580 -3980 -1520 -3920
rect -1480 -3980 -1420 -3920
rect -1380 -3980 -1320 -3920
rect -1280 -3980 -1220 -3920
rect -1180 -3980 -1120 -3920
rect -1080 -3980 -1020 -3920
rect -980 -3980 -920 -3920
rect -880 -3980 -820 -3920
rect -780 -3980 -720 -3920
rect -680 -3980 -620 -3920
rect -580 -3980 -520 -3920
rect -2380 -4080 -2320 -4020
rect -2280 -4080 -2220 -4020
rect -2180 -4080 -2120 -4020
rect -2080 -4080 -2020 -4020
rect -1980 -4080 -1920 -4020
rect -1880 -4080 -1820 -4020
rect -1780 -4080 -1720 -4020
rect -1680 -4080 -1620 -4020
rect -1580 -4080 -1520 -4020
rect -1480 -4080 -1420 -4020
rect -1380 -4080 -1320 -4020
rect -1280 -4080 -1220 -4020
rect -1180 -4080 -1120 -4020
rect -1080 -4080 -1020 -4020
rect -980 -4080 -920 -4020
rect -880 -4080 -820 -4020
rect -780 -4080 -720 -4020
rect -680 -4080 -620 -4020
rect -580 -4080 -520 -4020
<< metal1 >>
rect -2400 2080 -500 2100
rect -2400 2020 -2380 2080
rect -2320 2020 -2280 2080
rect -2220 2020 -2180 2080
rect -2120 2020 -2080 2080
rect -2020 2020 -1980 2080
rect -1920 2020 -1880 2080
rect -1820 2020 -1780 2080
rect -1720 2020 -1680 2080
rect -1620 2020 -1580 2080
rect -1520 2020 -1480 2080
rect -1420 2020 -1380 2080
rect -1320 2020 -1280 2080
rect -1220 2020 -1180 2080
rect -1120 2020 -1080 2080
rect -1020 2020 -980 2080
rect -920 2020 -880 2080
rect -820 2020 -780 2080
rect -720 2020 -680 2080
rect -620 2020 -580 2080
rect -520 2020 -500 2080
rect -2400 1980 -500 2020
rect -2400 1920 -2380 1980
rect -2320 1920 -2280 1980
rect -2220 1920 -2180 1980
rect -2120 1920 -2080 1980
rect -2020 1920 -1980 1980
rect -1920 1920 -1880 1980
rect -1820 1920 -1780 1980
rect -1720 1920 -1680 1980
rect -1620 1920 -1580 1980
rect -1520 1920 -1480 1980
rect -1420 1920 -1380 1980
rect -1320 1920 -1280 1980
rect -1220 1920 -1180 1980
rect -1120 1920 -1080 1980
rect -1020 1920 -980 1980
rect -920 1920 -880 1980
rect -820 1920 -780 1980
rect -720 1920 -680 1980
rect -620 1920 -580 1980
rect -520 1920 -500 1980
rect -2400 1880 -500 1920
rect -2400 1820 -2380 1880
rect -2320 1820 -2280 1880
rect -2220 1820 -2180 1880
rect -2120 1820 -2080 1880
rect -2020 1820 -1980 1880
rect -1920 1820 -1880 1880
rect -1820 1820 -1780 1880
rect -1720 1820 -1680 1880
rect -1620 1820 -1580 1880
rect -1520 1820 -1480 1880
rect -1420 1820 -1380 1880
rect -1320 1820 -1280 1880
rect -1220 1820 -1180 1880
rect -1120 1820 -1080 1880
rect -1020 1820 -980 1880
rect -920 1820 -880 1880
rect -820 1820 -780 1880
rect -720 1820 -680 1880
rect -620 1820 -580 1880
rect -520 1820 -500 1880
rect -2400 1780 -500 1820
rect -2400 1720 -2380 1780
rect -2320 1720 -2280 1780
rect -2220 1720 -2180 1780
rect -2120 1720 -2080 1780
rect -2020 1720 -1980 1780
rect -1920 1720 -1880 1780
rect -1820 1720 -1780 1780
rect -1720 1720 -1680 1780
rect -1620 1720 -1580 1780
rect -1520 1720 -1480 1780
rect -1420 1720 -1380 1780
rect -1320 1720 -1280 1780
rect -1220 1720 -1180 1780
rect -1120 1720 -1080 1780
rect -1020 1720 -980 1780
rect -920 1720 -880 1780
rect -820 1720 -780 1780
rect -720 1720 -680 1780
rect -620 1720 -580 1780
rect -520 1720 -500 1780
rect -2400 1680 -500 1720
rect -2400 1620 -2380 1680
rect -2320 1620 -2280 1680
rect -2220 1620 -2180 1680
rect -2120 1620 -2080 1680
rect -2020 1620 -1980 1680
rect -1920 1620 -1880 1680
rect -1820 1620 -1780 1680
rect -1720 1620 -1680 1680
rect -1620 1620 -1580 1680
rect -1520 1620 -1480 1680
rect -1420 1620 -1380 1680
rect -1320 1620 -1280 1680
rect -1220 1620 -1180 1680
rect -1120 1620 -1080 1680
rect -1020 1620 -980 1680
rect -920 1620 -880 1680
rect -820 1620 -780 1680
rect -720 1620 -680 1680
rect -620 1620 -580 1680
rect -520 1620 -500 1680
rect -2400 1580 -500 1620
rect -2400 1520 -2380 1580
rect -2320 1520 -2280 1580
rect -2220 1520 -2180 1580
rect -2120 1520 -2080 1580
rect -2020 1520 -1980 1580
rect -1920 1520 -1880 1580
rect -1820 1520 -1780 1580
rect -1720 1520 -1680 1580
rect -1620 1520 -1580 1580
rect -1520 1520 -1480 1580
rect -1420 1520 -1380 1580
rect -1320 1520 -1280 1580
rect -1220 1520 -1180 1580
rect -1120 1520 -1080 1580
rect -1020 1520 -980 1580
rect -920 1520 -880 1580
rect -820 1520 -780 1580
rect -720 1520 -680 1580
rect -620 1520 -580 1580
rect -520 1520 -500 1580
rect -2400 1480 -500 1520
rect -2400 1420 -2380 1480
rect -2320 1420 -2280 1480
rect -2220 1420 -2180 1480
rect -2120 1420 -2080 1480
rect -2020 1420 -1980 1480
rect -1920 1420 -1880 1480
rect -1820 1420 -1780 1480
rect -1720 1420 -1680 1480
rect -1620 1420 -1580 1480
rect -1520 1420 -1480 1480
rect -1420 1420 -1380 1480
rect -1320 1420 -1280 1480
rect -1220 1420 -1180 1480
rect -1120 1420 -1080 1480
rect -1020 1420 -980 1480
rect -920 1420 -880 1480
rect -820 1420 -780 1480
rect -720 1420 -680 1480
rect -620 1420 -580 1480
rect -520 1420 -500 1480
rect -2400 1400 -500 1420
rect -2180 880 -2080 900
rect -2180 820 -2160 880
rect -2100 820 -2080 880
rect -2180 780 -2080 820
rect -2180 720 -2160 780
rect -2100 720 -2080 780
rect -2180 700 -2080 720
rect -1560 880 -1460 900
rect -1560 820 -1540 880
rect -1480 820 -1460 880
rect -1560 780 -1460 820
rect -1560 720 -1540 780
rect -1480 720 -1460 780
rect -1560 700 -1460 720
rect -940 880 -840 900
rect -940 820 -920 880
rect -860 820 -840 880
rect -940 780 -840 820
rect -940 720 -920 780
rect -860 720 -840 780
rect -940 700 -840 720
rect -780 460 -680 1040
rect -180 460 -80 1040
rect 440 460 540 1040
rect -2200 360 540 460
rect 1200 500 1300 1100
rect 1780 880 1900 900
rect 1780 820 1800 880
rect 1860 820 1900 880
rect 1780 780 1900 820
rect 1780 720 1800 780
rect 1860 720 1900 780
rect 1780 700 1900 720
rect 2400 500 2500 1100
rect 3020 880 3140 900
rect 3020 820 3060 880
rect 3120 820 3140 880
rect 3020 780 3140 820
rect 3020 720 3060 780
rect 3120 720 3140 780
rect 3020 700 3140 720
rect 3600 500 3700 1100
rect 1200 400 3700 500
rect 4000 1000 5600 1200
rect 4000 880 4200 1000
rect 4000 820 4020 880
rect 4080 820 4120 880
rect 4180 820 4200 880
rect 4000 780 4200 820
rect 4000 720 4020 780
rect 4080 720 4120 780
rect 4180 720 4200 780
rect 1000 380 3900 400
rect -1940 -340 -1840 360
rect -2040 -400 -1840 -340
rect -1940 -440 -1840 -400
rect -2180 -620 -2080 -440
rect -1980 -620 -1840 -440
rect -2180 -900 -2100 -620
rect -1940 -660 -1840 -620
rect -2040 -720 -1840 -660
rect -1340 280 -1240 300
rect -1340 220 -1320 280
rect -1260 220 -1240 280
rect -1340 180 -1240 220
rect -1340 120 -1320 180
rect -1260 120 -1240 180
rect -1340 -900 -1240 120
rect -1176 -88 -436 -72
rect -2180 -940 -1240 -900
rect -1190 -182 -436 -88
rect -1190 -940 -1058 -182
rect -900 -920 -660 -240
rect -2180 -1000 -1000 -940
rect -1240 -1040 -1000 -1000
rect -1240 -1100 -1220 -1040
rect -1160 -1100 -1080 -1040
rect -1020 -1100 -1000 -1040
rect -1240 -1120 -1000 -1100
rect -1240 -1180 -1220 -1120
rect -1160 -1180 -1080 -1120
rect -1020 -1180 -1000 -1120
rect -1240 -1200 -1000 -1180
rect -2200 -2000 -1800 -1700
rect -900 -1780 -740 -920
rect -580 -940 -472 -182
rect -380 -920 -280 360
rect 1000 320 1020 380
rect 1080 320 1100 380
rect 1160 320 1180 380
rect 1240 320 3660 380
rect 3720 320 3740 380
rect 3800 320 3820 380
rect 3880 320 3900 380
rect 1000 280 3900 320
rect 1000 220 1020 280
rect 1080 220 1100 280
rect 1160 220 1180 280
rect 1240 220 1520 280
rect 1580 220 1920 280
rect 1980 220 2920 280
rect 2980 220 3320 280
rect 3380 220 3660 280
rect 3720 220 3740 280
rect 3800 220 3820 280
rect 3880 220 3900 280
rect 1000 200 3900 220
rect 4000 80 4200 720
rect 4340 580 4440 600
rect 4340 520 4360 580
rect 4420 520 4440 580
rect 4340 480 4440 520
rect 4340 420 4360 480
rect 4420 420 4440 480
rect 4340 400 4440 420
rect 4920 580 5020 600
rect 4920 520 4940 580
rect 5000 520 5020 580
rect 4920 480 5020 520
rect 4920 420 4940 480
rect 5000 420 5020 480
rect 4920 400 5020 420
rect 5540 580 5640 600
rect 5540 520 5560 580
rect 5620 520 5640 580
rect 5540 480 5640 520
rect 5540 420 5560 480
rect 5620 420 5640 480
rect 5540 400 5640 420
rect 4000 20 4020 80
rect 4080 20 4120 80
rect 4180 20 4200 80
rect 4000 0 4200 20
rect 4000 -20 5600 0
rect 4000 -80 4020 -20
rect 4080 -80 4120 -20
rect 4180 -80 5600 -20
rect 2410 -120 2490 -100
rect 2410 -180 2420 -120
rect 2480 -180 2490 -120
rect 2410 -220 2490 -180
rect 4000 -200 5600 -80
rect 2040 -240 2140 -220
rect 2040 -300 2060 -240
rect 2120 -300 2140 -240
rect 2040 -320 2140 -300
rect 2400 -280 2420 -220
rect 2480 -280 2500 -220
rect 2400 -320 2500 -280
rect 2740 -240 2840 -220
rect 2740 -300 2760 -240
rect 2820 -300 2840 -240
rect 2740 -320 2840 -300
rect 2410 -380 2420 -320
rect 2480 -380 2490 -320
rect 1440 -400 1600 -380
rect 1880 -400 2040 -380
rect 1440 -460 1520 -400
rect 1580 -460 1600 -400
rect 1440 -520 1600 -460
rect 1440 -580 1520 -520
rect 1580 -580 1600 -520
rect 1440 -600 1600 -580
rect 1700 -420 1800 -400
rect 1700 -480 1720 -420
rect 1780 -480 1800 -420
rect 1700 -500 1800 -480
rect 1700 -560 1720 -500
rect 1780 -560 1800 -500
rect 1700 -580 1800 -560
rect 1700 -640 1720 -580
rect 1780 -640 1800 -580
rect 1880 -460 1920 -400
rect 1980 -460 2040 -400
rect 1880 -520 2040 -460
rect 1880 -580 1920 -520
rect 1980 -580 2040 -520
rect 1880 -600 2040 -580
rect 2410 -420 2490 -380
rect 2410 -480 2420 -420
rect 2480 -480 2490 -420
rect 2410 -520 2490 -480
rect 2410 -580 2420 -520
rect 2480 -580 2490 -520
rect 1340 -800 1440 -640
rect 1700 -660 1800 -640
rect 1700 -720 1720 -660
rect 1780 -720 1800 -660
rect 1700 -740 1800 -720
rect 1700 -800 1720 -740
rect 1780 -800 1800 -740
rect 2410 -620 2490 -580
rect 2820 -400 2980 -380
rect 2820 -460 2900 -400
rect 2960 -460 2980 -400
rect 2820 -520 2980 -460
rect 2820 -580 2900 -520
rect 2960 -580 2980 -520
rect 2820 -600 2980 -580
rect 3300 -400 3460 -380
rect 3300 -460 3320 -400
rect 3380 -460 3460 -400
rect 3300 -520 3460 -460
rect 3300 -580 3320 -520
rect 3380 -580 3460 -520
rect 3300 -600 3460 -580
rect 2410 -680 2420 -620
rect 2480 -680 2490 -620
rect 2410 -700 2490 -680
rect 2410 -760 2420 -700
rect 2480 -760 2490 -700
rect 3440 -800 3540 -640
rect 100 -820 3900 -800
rect 100 -880 1720 -820
rect 1780 -880 3900 -820
rect 100 -900 3900 -880
rect -640 -1040 -400 -940
rect -640 -1100 -620 -1040
rect -560 -1100 -480 -1040
rect -420 -1100 -400 -1040
rect -640 -1120 -400 -1100
rect -640 -1180 -620 -1120
rect -560 -1180 -480 -1120
rect -420 -1180 -400 -1120
rect -640 -1200 -400 -1180
rect -820 -1820 -720 -1780
rect -1100 -2400 -700 -2100
rect -2200 -2700 -1800 -2400
rect -2200 -3400 -1780 -2900
rect -1100 -3000 -700 -2700
rect -2400 -3420 -500 -3400
rect -2400 -3480 -2380 -3420
rect -2320 -3480 -2280 -3420
rect -2220 -3480 -2180 -3420
rect -2120 -3480 -2080 -3420
rect -2020 -3480 -1980 -3420
rect -1920 -3480 -1880 -3420
rect -1820 -3480 -1780 -3420
rect -1720 -3480 -1680 -3420
rect -1620 -3480 -1580 -3420
rect -1520 -3480 -1480 -3420
rect -1420 -3480 -1380 -3420
rect -1320 -3480 -1280 -3420
rect -1220 -3480 -1180 -3420
rect -1120 -3480 -1080 -3420
rect -1020 -3480 -980 -3420
rect -920 -3480 -880 -3420
rect -820 -3480 -780 -3420
rect -720 -3480 -680 -3420
rect -620 -3480 -580 -3420
rect -520 -3480 -500 -3420
rect -2400 -3520 -500 -3480
rect -2400 -3580 -2380 -3520
rect -2320 -3580 -2280 -3520
rect -2220 -3580 -2180 -3520
rect -2120 -3580 -2080 -3520
rect -2020 -3580 -1980 -3520
rect -1920 -3580 -1880 -3520
rect -1820 -3580 -1780 -3520
rect -1720 -3580 -1680 -3520
rect -1620 -3580 -1580 -3520
rect -1520 -3580 -1480 -3520
rect -1420 -3580 -1380 -3520
rect -1320 -3580 -1280 -3520
rect -1220 -3580 -1180 -3520
rect -1120 -3580 -1080 -3520
rect -1020 -3580 -980 -3520
rect -920 -3580 -880 -3520
rect -820 -3580 -780 -3520
rect -720 -3580 -680 -3520
rect -620 -3580 -580 -3520
rect -520 -3580 -500 -3520
rect -2400 -3620 -500 -3580
rect -2400 -3680 -2380 -3620
rect -2320 -3680 -2280 -3620
rect -2220 -3680 -2180 -3620
rect -2120 -3680 -2080 -3620
rect -2020 -3680 -1980 -3620
rect -1920 -3680 -1880 -3620
rect -1820 -3680 -1780 -3620
rect -1720 -3680 -1680 -3620
rect -1620 -3680 -1580 -3620
rect -1520 -3680 -1480 -3620
rect -1420 -3680 -1380 -3620
rect -1320 -3680 -1280 -3620
rect -1220 -3680 -1180 -3620
rect -1120 -3680 -1080 -3620
rect -1020 -3680 -980 -3620
rect -920 -3680 -880 -3620
rect -820 -3680 -780 -3620
rect -720 -3680 -680 -3620
rect -620 -3680 -580 -3620
rect -520 -3680 -500 -3620
rect -2400 -3720 -500 -3680
rect -2400 -3780 -2380 -3720
rect -2320 -3780 -2280 -3720
rect -2220 -3780 -2180 -3720
rect -2120 -3780 -2080 -3720
rect -2020 -3780 -1980 -3720
rect -1920 -3780 -1880 -3720
rect -1820 -3780 -1780 -3720
rect -1720 -3780 -1680 -3720
rect -1620 -3780 -1580 -3720
rect -1520 -3780 -1480 -3720
rect -1420 -3780 -1380 -3720
rect -1320 -3780 -1280 -3720
rect -1220 -3780 -1180 -3720
rect -1120 -3780 -1080 -3720
rect -1020 -3780 -980 -3720
rect -920 -3780 -880 -3720
rect -820 -3780 -780 -3720
rect -720 -3780 -680 -3720
rect -620 -3780 -580 -3720
rect -520 -3780 -500 -3720
rect -2400 -3820 -500 -3780
rect -2400 -3880 -2380 -3820
rect -2320 -3880 -2280 -3820
rect -2220 -3880 -2180 -3820
rect -2120 -3880 -2080 -3820
rect -2020 -3880 -1980 -3820
rect -1920 -3880 -1880 -3820
rect -1820 -3880 -1780 -3820
rect -1720 -3880 -1680 -3820
rect -1620 -3880 -1580 -3820
rect -1520 -3880 -1480 -3820
rect -1420 -3880 -1380 -3820
rect -1320 -3880 -1280 -3820
rect -1220 -3880 -1180 -3820
rect -1120 -3880 -1080 -3820
rect -1020 -3880 -980 -3820
rect -920 -3880 -880 -3820
rect -820 -3880 -780 -3820
rect -720 -3880 -680 -3820
rect -620 -3880 -580 -3820
rect -520 -3880 -500 -3820
rect -2400 -3920 -500 -3880
rect -2400 -3980 -2380 -3920
rect -2320 -3980 -2280 -3920
rect -2220 -3980 -2180 -3920
rect -2120 -3980 -2080 -3920
rect -2020 -3980 -1980 -3920
rect -1920 -3980 -1880 -3920
rect -1820 -3980 -1780 -3920
rect -1720 -3980 -1680 -3920
rect -1620 -3980 -1580 -3920
rect -1520 -3980 -1480 -3920
rect -1420 -3980 -1380 -3920
rect -1320 -3980 -1280 -3920
rect -1220 -3980 -1180 -3920
rect -1120 -3980 -1080 -3920
rect -1020 -3980 -980 -3920
rect -920 -3980 -880 -3920
rect -820 -3980 -780 -3920
rect -720 -3980 -680 -3920
rect -620 -3980 -580 -3920
rect -520 -3980 -500 -3920
rect -2400 -4020 -500 -3980
rect -2400 -4080 -2380 -4020
rect -2320 -4080 -2280 -4020
rect -2220 -4080 -2180 -4020
rect -2120 -4080 -2080 -4020
rect -2020 -4080 -1980 -4020
rect -1920 -4080 -1880 -4020
rect -1820 -4080 -1780 -4020
rect -1720 -4080 -1680 -4020
rect -1620 -4080 -1580 -4020
rect -1520 -4080 -1480 -4020
rect -1420 -4080 -1380 -4020
rect -1320 -4080 -1280 -4020
rect -1220 -4080 -1180 -4020
rect -1120 -4080 -1080 -4020
rect -1020 -4080 -980 -4020
rect -920 -4080 -880 -4020
rect -820 -4080 -780 -4020
rect -720 -4080 -680 -4020
rect -620 -4080 -580 -4020
rect -520 -4080 -500 -4020
rect -2400 -4100 -500 -4080
rect 100 -4380 200 -900
rect 3100 -1000 3120 -980
rect 400 -1040 3120 -1000
rect 3180 -1000 3200 -980
rect 3180 -1040 3900 -1000
rect 400 -1060 3900 -1040
rect 400 -1100 3120 -1060
rect 400 -4380 500 -1100
rect 1340 -1240 1440 -1100
rect 3100 -1120 3120 -1100
rect 3180 -1100 3900 -1060
rect 3180 -1120 3200 -1100
rect 3100 -1140 3200 -1120
rect 2410 -1200 2420 -1140
rect 2480 -1200 2490 -1140
rect 2410 -1220 2490 -1200
rect 2410 -1280 2420 -1220
rect 2480 -1280 2490 -1220
rect 3100 -1200 3120 -1140
rect 3180 -1200 3200 -1140
rect 3100 -1220 3200 -1200
rect 3100 -1280 3120 -1220
rect 3180 -1280 3200 -1220
rect 3440 -1240 3540 -1100
rect 1200 -1300 1360 -1280
rect 1200 -1360 1220 -1300
rect 1280 -1360 1360 -1300
rect 1200 -1420 1360 -1360
rect 1200 -1480 1220 -1420
rect 1280 -1480 1360 -1420
rect 1200 -1500 1360 -1480
rect 1900 -1300 2060 -1280
rect 1900 -1360 1920 -1300
rect 1980 -1360 2060 -1300
rect 1900 -1420 2060 -1360
rect 1900 -1480 1920 -1420
rect 1980 -1480 2060 -1420
rect 1900 -1500 2060 -1480
rect 2410 -1320 2490 -1280
rect 2410 -1380 2420 -1320
rect 2480 -1380 2490 -1320
rect 2410 -1420 2490 -1380
rect 2410 -1480 2420 -1420
rect 2480 -1480 2490 -1420
rect 2410 -1520 2490 -1480
rect 2820 -1300 3000 -1280
rect 2820 -1360 2920 -1300
rect 2980 -1360 3000 -1300
rect 2820 -1420 3000 -1360
rect 2820 -1480 2920 -1420
rect 2980 -1480 3000 -1420
rect 3100 -1300 3200 -1280
rect 3100 -1360 3120 -1300
rect 3180 -1360 3200 -1300
rect 3100 -1380 3200 -1360
rect 3100 -1440 3120 -1380
rect 3180 -1440 3200 -1380
rect 3100 -1460 3200 -1440
rect 3520 -1300 3680 -1280
rect 3520 -1360 3560 -1300
rect 3620 -1360 3680 -1300
rect 3520 -1420 3680 -1360
rect 2820 -1500 3000 -1480
rect 3520 -1480 3560 -1420
rect 3620 -1480 3680 -1420
rect 3520 -1500 3680 -1480
rect 4000 -1300 4200 -200
rect 4340 -700 4440 -680
rect 4340 -760 4360 -700
rect 4420 -760 4440 -700
rect 4340 -800 4440 -760
rect 4340 -860 4360 -800
rect 4420 -860 4440 -800
rect 4340 -880 4440 -860
rect 4940 -700 5040 -680
rect 4940 -760 4960 -700
rect 5020 -760 5040 -700
rect 4940 -800 5040 -760
rect 4940 -860 4960 -800
rect 5020 -860 5040 -800
rect 4940 -880 5040 -860
rect 5540 -700 5640 -680
rect 5540 -760 5560 -700
rect 5620 -760 5640 -700
rect 5540 -800 5640 -760
rect 5540 -860 5560 -800
rect 5620 -860 5640 -800
rect 5540 -880 5640 -860
rect 4000 -1500 5600 -1300
rect 2410 -1540 2420 -1520
rect 2040 -1560 2140 -1540
rect 2040 -1620 2060 -1560
rect 2120 -1620 2140 -1560
rect 2040 -1640 2140 -1620
rect 2400 -1580 2420 -1540
rect 2480 -1540 2490 -1520
rect 2480 -1580 2500 -1540
rect 2400 -1620 2500 -1580
rect 2400 -1640 2420 -1620
rect 2410 -1680 2420 -1640
rect 2480 -1640 2500 -1620
rect 2740 -1560 2840 -1540
rect 2740 -1620 2760 -1560
rect 2820 -1620 2840 -1560
rect 2740 -1640 2840 -1620
rect 2480 -1680 2490 -1640
rect 2410 -1700 2490 -1680
rect 2400 -1720 2500 -1700
rect 2400 -1780 2420 -1720
rect 2480 -1780 2500 -1720
rect 2400 -2000 2500 -1780
rect 1940 -2080 2500 -2000
rect 4000 -1820 4200 -1500
rect 4000 -1880 4020 -1820
rect 4080 -1880 4120 -1820
rect 4180 -1880 4200 -1820
rect 4000 -1920 4200 -1880
rect 4000 -1980 4020 -1920
rect 4080 -1980 4120 -1920
rect 4180 -1980 4200 -1920
rect 1160 -2120 1400 -2100
rect 1160 -2180 1180 -2120
rect 1240 -2180 1320 -2120
rect 1380 -2180 1400 -2120
rect 1160 -2220 1400 -2180
rect 1160 -2280 1180 -2220
rect 1240 -2280 1320 -2220
rect 1380 -2280 1400 -2220
rect 1160 -2360 1400 -2280
rect 1420 -3200 1520 -2400
rect 1940 -3200 2040 -2080
rect 2560 -2140 2800 -2120
rect 2560 -2200 2580 -2140
rect 2640 -2200 2720 -2140
rect 2780 -2200 2800 -2140
rect 2560 -2220 2800 -2200
rect 2560 -2280 2580 -2220
rect 2640 -2280 2720 -2220
rect 2780 -2280 2800 -2220
rect 2560 -2440 2800 -2280
rect 2880 -2140 3120 -2120
rect 2880 -2200 2900 -2140
rect 2960 -2200 3040 -2140
rect 3100 -2200 3120 -2140
rect 2880 -2220 3120 -2200
rect 2880 -2280 2900 -2220
rect 2960 -2280 3040 -2220
rect 3100 -2280 3120 -2220
rect 2880 -2440 3120 -2280
rect 3180 -2140 3420 -2120
rect 3180 -2200 3200 -2140
rect 3260 -2200 3340 -2140
rect 3400 -2200 3420 -2140
rect 3180 -2220 3420 -2200
rect 3180 -2280 3200 -2220
rect 3260 -2280 3340 -2220
rect 3400 -2280 3420 -2220
rect 3180 -2440 3420 -2280
rect 3480 -2140 3720 -2120
rect 3480 -2200 3500 -2140
rect 3560 -2200 3640 -2140
rect 3700 -2200 3720 -2140
rect 3480 -2220 3720 -2200
rect 3480 -2280 3500 -2220
rect 3560 -2280 3640 -2220
rect 3700 -2280 3720 -2220
rect 3480 -2440 3720 -2280
rect 4000 -2600 4200 -1980
rect 4340 -1980 4440 -1960
rect 4340 -2040 4360 -1980
rect 4420 -2040 4440 -1980
rect 4340 -2080 4440 -2040
rect 4340 -2140 4360 -2080
rect 4420 -2140 4440 -2080
rect 4340 -2160 4440 -2140
rect 4940 -1980 5040 -1960
rect 4940 -2040 4960 -1980
rect 5020 -2040 5040 -1980
rect 4940 -2080 5040 -2040
rect 4940 -2140 4960 -2080
rect 5020 -2140 5040 -2080
rect 4940 -2160 5040 -2140
rect 5540 -1980 5640 -1960
rect 5540 -2040 5560 -1980
rect 5620 -2040 5640 -1980
rect 5540 -2080 5640 -2040
rect 5540 -2140 5560 -2080
rect 5620 -2140 5640 -2080
rect 5540 -2160 5640 -2140
rect 2500 -2720 2600 -2700
rect 2500 -2780 2520 -2720
rect 2580 -2780 2600 -2720
rect 2500 -2820 2600 -2780
rect 2500 -2880 2520 -2820
rect 2580 -2880 2600 -2820
rect 2500 -2900 2600 -2880
rect 3100 -2720 3200 -2700
rect 3100 -2780 3120 -2720
rect 3180 -2780 3200 -2720
rect 3100 -2820 3200 -2780
rect 3100 -2880 3120 -2820
rect 3180 -2880 3200 -2820
rect 3100 -2900 3200 -2880
rect 3720 -2720 3820 -2700
rect 3720 -2780 3740 -2720
rect 3800 -2780 3820 -2720
rect 3720 -2820 3820 -2780
rect 3720 -2880 3740 -2820
rect 3800 -2880 3820 -2820
rect 3720 -2900 3820 -2880
rect 4000 -2800 5600 -2600
rect 1420 -3300 2040 -3200
rect 4000 -3800 4200 -2800
rect 4340 -3260 4440 -3240
rect 4340 -3320 4360 -3260
rect 4420 -3320 4440 -3260
rect 4340 -3360 4440 -3320
rect 4340 -3420 4360 -3360
rect 4420 -3420 4440 -3360
rect 4340 -3440 4440 -3420
rect 4920 -3260 5020 -3240
rect 4920 -3320 4940 -3260
rect 5000 -3320 5020 -3260
rect 4920 -3360 5020 -3320
rect 4920 -3420 4940 -3360
rect 5000 -3420 5020 -3360
rect 4920 -3440 5020 -3420
rect 5540 -3260 5640 -3240
rect 5540 -3320 5560 -3260
rect 5620 -3320 5640 -3260
rect 5540 -3360 5640 -3320
rect 5540 -3420 5560 -3360
rect 5620 -3420 5640 -3360
rect 5540 -3440 5640 -3420
rect 4000 -4000 5600 -3800
rect 40 -4580 240 -4380
rect 360 -4580 560 -4380
rect 4340 -4520 4440 -4500
rect 4340 -4580 4360 -4520
rect 4420 -4580 4440 -4520
rect 4340 -4620 4440 -4580
rect 4340 -4680 4360 -4620
rect 4420 -4680 4440 -4620
rect 4340 -4700 4440 -4680
rect 4920 -4520 5020 -4500
rect 4920 -4580 4940 -4520
rect 5000 -4580 5020 -4520
rect 4920 -4620 5020 -4580
rect 4920 -4680 4940 -4620
rect 5000 -4680 5020 -4620
rect 4920 -4700 5020 -4680
rect 5540 -4520 5640 -4500
rect 5540 -4580 5560 -4520
rect 5620 -4580 5640 -4520
rect 5540 -4620 5640 -4580
rect 5540 -4680 5560 -4620
rect 5620 -4680 5640 -4620
rect 5540 -4700 5640 -4680
rect 3700 -5120 3900 -5100
rect 3700 -5180 3720 -5120
rect 3780 -5180 3820 -5120
rect 3880 -5180 3900 -5120
rect 3700 -5220 3900 -5180
rect 3700 -5280 3720 -5220
rect 3780 -5280 3820 -5220
rect 3880 -5280 3900 -5220
rect 3700 -5300 3900 -5280
<< via1 >>
rect -2160 820 -2100 880
rect -2160 720 -2100 780
rect -1540 820 -1480 880
rect -1540 720 -1480 780
rect -920 820 -860 880
rect -920 720 -860 780
rect 1800 820 1860 880
rect 1800 720 1860 780
rect 3060 820 3120 880
rect 3060 720 3120 780
rect 4020 820 4080 880
rect 4120 820 4180 880
rect 4020 720 4080 780
rect 4120 720 4180 780
rect -1320 220 -1260 280
rect -1320 120 -1260 180
rect -1220 -1100 -1160 -1040
rect -1080 -1100 -1020 -1040
rect -1220 -1180 -1160 -1120
rect -1080 -1180 -1020 -1120
rect 1020 320 1080 380
rect 1100 320 1160 380
rect 1180 320 1240 380
rect 3660 320 3720 380
rect 3740 320 3800 380
rect 3820 320 3880 380
rect 1020 220 1080 280
rect 1100 220 1160 280
rect 1180 220 1240 280
rect 1520 220 1580 280
rect 1920 220 1980 280
rect 2920 220 2980 280
rect 3320 220 3380 280
rect 3660 220 3720 280
rect 3740 220 3800 280
rect 3820 220 3880 280
rect 4360 520 4420 580
rect 4360 420 4420 480
rect 4940 520 5000 580
rect 4940 420 5000 480
rect 5560 520 5620 580
rect 5560 420 5620 480
rect 4020 20 4080 80
rect 4120 20 4180 80
rect 4020 -80 4080 -20
rect 4120 -80 4180 -20
rect 2060 -300 2120 -240
rect 2760 -300 2820 -240
rect 1520 -460 1580 -400
rect 1520 -580 1580 -520
rect 1720 -480 1780 -420
rect 1720 -560 1780 -500
rect 1720 -640 1780 -580
rect 1920 -460 1980 -400
rect 1920 -580 1980 -520
rect 1720 -720 1780 -660
rect 1720 -800 1780 -740
rect 2900 -460 2960 -400
rect 2900 -580 2960 -520
rect 3320 -460 3380 -400
rect 3320 -580 3380 -520
rect 2420 -760 2480 -700
rect 1720 -880 1780 -820
rect -620 -1100 -560 -1040
rect -480 -1100 -420 -1040
rect -620 -1180 -560 -1120
rect -480 -1180 -420 -1120
rect 3120 -1040 3180 -980
rect 3120 -1120 3180 -1060
rect 2420 -1200 2480 -1140
rect 3120 -1200 3180 -1140
rect 3120 -1280 3180 -1220
rect 1220 -1360 1280 -1300
rect 1220 -1480 1280 -1420
rect 1920 -1360 1980 -1300
rect 1920 -1480 1980 -1420
rect 2920 -1360 2980 -1300
rect 2920 -1480 2980 -1420
rect 3120 -1360 3180 -1300
rect 3120 -1440 3180 -1380
rect 3560 -1360 3620 -1300
rect 3560 -1480 3620 -1420
rect 4360 -760 4420 -700
rect 4360 -860 4420 -800
rect 4960 -760 5020 -700
rect 4960 -860 5020 -800
rect 5560 -760 5620 -700
rect 5560 -860 5620 -800
rect 2060 -1620 2120 -1560
rect 2760 -1620 2820 -1560
rect 4020 -1880 4080 -1820
rect 4120 -1880 4180 -1820
rect 4020 -1980 4080 -1920
rect 4120 -1980 4180 -1920
rect 1180 -2180 1240 -2120
rect 1320 -2180 1380 -2120
rect 1180 -2280 1240 -2220
rect 1320 -2280 1380 -2220
rect 2580 -2200 2640 -2140
rect 2720 -2200 2780 -2140
rect 2580 -2280 2640 -2220
rect 2720 -2280 2780 -2220
rect 2900 -2200 2960 -2140
rect 3040 -2200 3100 -2140
rect 2900 -2280 2960 -2220
rect 3040 -2280 3100 -2220
rect 3200 -2200 3260 -2140
rect 3340 -2200 3400 -2140
rect 3200 -2280 3260 -2220
rect 3340 -2280 3400 -2220
rect 3500 -2200 3560 -2140
rect 3640 -2200 3700 -2140
rect 3500 -2280 3560 -2220
rect 3640 -2280 3700 -2220
rect 4360 -2040 4420 -1980
rect 4360 -2140 4420 -2080
rect 4960 -2040 5020 -1980
rect 4960 -2140 5020 -2080
rect 5560 -2040 5620 -1980
rect 5560 -2140 5620 -2080
rect 2520 -2780 2580 -2720
rect 2520 -2880 2580 -2820
rect 3120 -2780 3180 -2720
rect 3120 -2880 3180 -2820
rect 3740 -2780 3800 -2720
rect 3740 -2880 3800 -2820
rect 4360 -3320 4420 -3260
rect 4360 -3420 4420 -3360
rect 4940 -3320 5000 -3260
rect 4940 -3420 5000 -3360
rect 5560 -3320 5620 -3260
rect 5560 -3420 5620 -3360
rect 4360 -4580 4420 -4520
rect 4360 -4680 4420 -4620
rect 4940 -4580 5000 -4520
rect 4940 -4680 5000 -4620
rect 5560 -4580 5620 -4520
rect 5560 -4680 5620 -4620
rect 3720 -5180 3780 -5120
rect 3820 -5180 3880 -5120
rect 3720 -5280 3780 -5220
rect 3820 -5280 3880 -5220
<< metal2 >>
rect -2300 880 -800 900
rect -2300 820 -2160 880
rect -2100 820 -1540 880
rect -1480 820 -920 880
rect -860 820 -800 880
rect -2300 780 -800 820
rect -2300 720 -2160 780
rect -2100 720 -1540 780
rect -1480 720 -920 780
rect -860 720 -800 780
rect -2300 700 -800 720
rect 1100 880 4200 900
rect 1100 820 1800 880
rect 1860 820 3060 880
rect 3120 820 4020 880
rect 4080 820 4120 880
rect 4180 820 4200 880
rect 1100 780 4200 820
rect 1100 720 1800 780
rect 1860 720 3060 780
rect 3120 720 4020 780
rect 4080 720 4120 780
rect 4180 720 4200 780
rect 1100 700 4200 720
rect -1600 300 -1440 700
rect 4340 580 5900 600
rect 4340 520 4360 580
rect 4420 520 4940 580
rect 5000 520 5560 580
rect 5620 520 5900 580
rect 4340 480 5900 520
rect 4340 420 4360 480
rect 4420 420 4940 480
rect 5000 420 5560 480
rect 5620 420 5900 480
rect 4340 400 5900 420
rect 1000 380 3900 400
rect 1000 320 1020 380
rect 1080 320 1100 380
rect 1160 320 1180 380
rect 1240 320 3660 380
rect 3720 320 3740 380
rect 3800 320 3820 380
rect 3880 320 3900 380
rect -2100 280 500 300
rect -2100 220 -1320 280
rect -1260 220 500 280
rect -2100 180 500 220
rect 1000 280 3900 320
rect 1000 220 1020 280
rect 1080 220 1100 280
rect 1160 220 1180 280
rect 1240 220 1520 280
rect 1580 220 1920 280
rect 1980 220 2920 280
rect 2980 220 3320 280
rect 3380 220 3660 280
rect 3720 220 3740 280
rect 3800 220 3820 280
rect 3880 220 3900 280
rect 1000 200 3900 220
rect -2100 120 -1320 180
rect -1260 120 500 180
rect -2100 100 500 120
rect 1100 80 4200 100
rect 1100 20 4020 80
rect 4080 20 4120 80
rect 4180 20 4200 80
rect 1100 -20 4200 20
rect 1100 -80 4020 -20
rect 4080 -80 4120 -20
rect 4180 -80 4200 -20
rect 1100 -100 4200 -80
rect -1300 -1040 0 -1000
rect -1300 -1100 -1220 -1040
rect -1160 -1100 -1080 -1040
rect -1020 -1100 -620 -1040
rect -560 -1100 -480 -1040
rect -420 -1100 0 -1040
rect -1300 -1120 0 -1100
rect -1300 -1180 -1220 -1120
rect -1160 -1180 -1080 -1120
rect -1020 -1180 -620 -1120
rect -560 -1180 -480 -1120
rect -420 -1180 0 -1120
rect -1300 -1200 0 -1180
rect -200 -2100 0 -1200
rect 1200 -1280 1300 -200
rect 1860 -380 1960 -100
rect 2000 -240 3200 -220
rect 2000 -300 2060 -240
rect 2120 -300 2760 -240
rect 2820 -300 3200 -240
rect 2000 -320 3200 -300
rect 1440 -400 1600 -380
rect 1860 -400 2040 -380
rect 1440 -460 1520 -400
rect 1580 -460 1600 -400
rect 1440 -520 1600 -460
rect 1440 -580 1520 -520
rect 1580 -580 1600 -520
rect 1440 -600 1600 -580
rect 1700 -420 1800 -400
rect 1700 -480 1720 -420
rect 1780 -480 1800 -420
rect 1700 -500 1800 -480
rect 1700 -560 1720 -500
rect 1780 -560 1800 -500
rect 1700 -580 1800 -560
rect 1700 -640 1720 -580
rect 1780 -640 1800 -580
rect 1700 -660 1800 -640
rect 1700 -720 1720 -660
rect 1780 -720 1800 -660
rect 1700 -740 1800 -720
rect 1700 -800 1720 -740
rect 1780 -800 1800 -740
rect 1860 -460 1920 -400
rect 1980 -440 2040 -400
rect 2820 -400 2980 -380
rect 2820 -440 2900 -400
rect 1980 -460 2900 -440
rect 2960 -460 2980 -400
rect 1860 -520 2980 -460
rect 1860 -580 1920 -520
rect 1980 -540 2900 -520
rect 1980 -580 2040 -540
rect 1860 -600 2040 -580
rect 2820 -580 2900 -540
rect 2960 -580 2980 -520
rect 2820 -600 2980 -580
rect 1860 -800 1960 -600
rect 2410 -700 2490 -690
rect 2410 -760 2420 -700
rect 2480 -760 2490 -700
rect 1700 -820 1800 -800
rect 1700 -880 1720 -820
rect 1780 -880 1800 -820
rect 1200 -1300 1360 -1280
rect 1200 -1360 1220 -1300
rect 1280 -1360 1360 -1300
rect 1200 -1420 1360 -1360
rect 1200 -1480 1220 -1420
rect 1280 -1480 1360 -1420
rect 1200 -1500 1360 -1480
rect 1200 -1800 1300 -1500
rect 1700 -1540 1800 -880
rect 2410 -1140 2490 -760
rect 2410 -1200 2420 -1140
rect 2480 -1200 2490 -1140
rect 2410 -1210 2490 -1200
rect 3100 -980 3200 -320
rect 3300 -400 3460 -380
rect 3300 -460 3320 -400
rect 3380 -460 3460 -400
rect 3300 -520 3460 -460
rect 3300 -580 3320 -520
rect 3380 -580 3460 -520
rect 3300 -600 3460 -580
rect 3100 -1040 3120 -980
rect 3180 -1040 3200 -980
rect 3100 -1060 3200 -1040
rect 3100 -1120 3120 -1060
rect 3180 -1120 3200 -1060
rect 3100 -1140 3200 -1120
rect 3100 -1200 3120 -1140
rect 3180 -1200 3200 -1140
rect 3100 -1220 3200 -1200
rect 3100 -1280 3120 -1220
rect 3180 -1280 3200 -1220
rect 3600 -1280 3700 -200
rect 5720 -680 5900 400
rect 4340 -700 5900 -680
rect 4340 -760 4360 -700
rect 4420 -760 4960 -700
rect 5020 -760 5560 -700
rect 5620 -760 5900 -700
rect 4340 -800 5900 -760
rect 4340 -860 4360 -800
rect 4420 -860 4960 -800
rect 5020 -860 5560 -800
rect 5620 -860 5900 -800
rect 4340 -880 5900 -860
rect 1900 -1300 2060 -1280
rect 1900 -1360 1920 -1300
rect 1980 -1360 2060 -1300
rect 1900 -1420 2060 -1360
rect 1900 -1480 1920 -1420
rect 1980 -1480 2060 -1420
rect 1900 -1500 2060 -1480
rect 2820 -1300 3000 -1280
rect 2820 -1360 2920 -1300
rect 2980 -1360 3000 -1300
rect 2820 -1420 3000 -1360
rect 2820 -1480 2920 -1420
rect 2980 -1480 3000 -1420
rect 3100 -1300 3200 -1280
rect 3100 -1360 3120 -1300
rect 3180 -1360 3200 -1300
rect 3100 -1380 3200 -1360
rect 3100 -1440 3120 -1380
rect 3180 -1440 3200 -1380
rect 3100 -1460 3200 -1440
rect 3520 -1300 3700 -1280
rect 3520 -1360 3560 -1300
rect 3620 -1360 3700 -1300
rect 3520 -1420 3700 -1360
rect 2820 -1500 3000 -1480
rect 3520 -1480 3560 -1420
rect 3620 -1480 3700 -1420
rect 3520 -1500 3700 -1480
rect 1700 -1560 2900 -1540
rect 1700 -1620 2060 -1560
rect 2120 -1620 2760 -1560
rect 2820 -1620 2900 -1560
rect 1700 -1640 2900 -1620
rect 3600 -1800 3700 -1500
rect 1100 -1820 4200 -1800
rect 1100 -1880 4020 -1820
rect 4080 -1880 4120 -1820
rect 4180 -1880 4200 -1820
rect 1100 -1920 4200 -1880
rect 1100 -1980 4020 -1920
rect 4080 -1980 4120 -1920
rect 4180 -1980 4200 -1920
rect 5720 -1960 5900 -880
rect 1100 -2000 4200 -1980
rect 4340 -1980 5900 -1960
rect 4340 -2040 4360 -1980
rect 4420 -2040 4960 -1980
rect 5020 -2040 5560 -1980
rect 5620 -2040 5900 -1980
rect 4340 -2080 5900 -2040
rect -200 -2120 3900 -2100
rect -200 -2180 1180 -2120
rect 1240 -2180 1320 -2120
rect 1380 -2140 3900 -2120
rect 1380 -2180 2580 -2140
rect -200 -2200 2580 -2180
rect 2640 -2200 2720 -2140
rect 2780 -2200 2900 -2140
rect 2960 -2200 3040 -2140
rect 3100 -2200 3200 -2140
rect 3260 -2200 3340 -2140
rect 3400 -2200 3500 -2140
rect 3560 -2200 3640 -2140
rect 3700 -2200 3900 -2140
rect 4340 -2140 4360 -2080
rect 4420 -2140 4960 -2080
rect 5020 -2140 5560 -2080
rect 5620 -2140 5900 -2080
rect 4340 -2160 5900 -2140
rect -200 -2220 3900 -2200
rect -200 -2280 1180 -2220
rect 1240 -2280 1320 -2220
rect 1380 -2280 2580 -2220
rect 2640 -2280 2720 -2220
rect 2780 -2280 2900 -2220
rect 2960 -2280 3040 -2220
rect 3100 -2280 3200 -2220
rect 3260 -2280 3340 -2220
rect 3400 -2280 3500 -2220
rect 3560 -2280 3640 -2220
rect 3700 -2280 3900 -2220
rect -200 -2300 3900 -2280
rect 5720 -2700 5900 -2160
rect 2500 -2720 5900 -2700
rect 2500 -2780 2520 -2720
rect 2580 -2780 3120 -2720
rect 3180 -2780 3740 -2720
rect 3800 -2780 5900 -2720
rect 2500 -2820 5900 -2780
rect 2500 -2880 2520 -2820
rect 2580 -2880 3120 -2820
rect 3180 -2880 3740 -2820
rect 3800 -2880 5900 -2820
rect 2500 -2900 5900 -2880
rect 5720 -3240 5900 -2900
rect 4340 -3260 5900 -3240
rect 4340 -3320 4360 -3260
rect 4420 -3320 4940 -3260
rect 5000 -3320 5560 -3260
rect 5620 -3320 5900 -3260
rect 4340 -3360 5900 -3320
rect 4340 -3420 4360 -3360
rect 4420 -3420 4940 -3360
rect 5000 -3420 5560 -3360
rect 5620 -3420 5900 -3360
rect 4340 -3440 5900 -3420
rect 5720 -4500 5900 -3440
rect 4340 -4520 5900 -4500
rect 4340 -4580 4360 -4520
rect 4420 -4580 4940 -4520
rect 5000 -4580 5560 -4520
rect 5620 -4580 5900 -4520
rect 4340 -4620 5900 -4580
rect 4340 -4680 4360 -4620
rect 4420 -4680 4940 -4620
rect 5000 -4680 5560 -4620
rect 5620 -4680 5900 -4620
rect 4340 -4700 5900 -4680
rect 5720 -5100 5900 -4700
rect 3700 -5120 5900 -5100
rect 3700 -5180 3720 -5120
rect 3780 -5180 3820 -5120
rect 3880 -5180 5640 -5120
rect 5700 -5180 5740 -5120
rect 5800 -5180 5900 -5120
rect 3700 -5220 5900 -5180
rect 3700 -5280 3720 -5220
rect 3780 -5280 3820 -5220
rect 3880 -5280 5640 -5220
rect 5700 -5280 5740 -5220
rect 5800 -5280 5900 -5220
rect 3700 -5300 5900 -5280
<< via2 >>
rect 4020 820 4080 880
rect 4120 820 4180 880
rect 4020 720 4080 780
rect 4120 720 4180 780
rect 1520 220 1580 280
rect 1920 220 1980 280
rect 2920 220 2980 280
rect 3320 220 3380 280
rect 1520 -460 1580 -400
rect 1520 -580 1580 -520
rect 3320 -460 3380 -400
rect 3320 -580 3380 -520
rect 1920 -1360 1980 -1300
rect 1920 -1480 1980 -1420
rect 2920 -1360 2980 -1300
rect 2920 -1480 2980 -1420
rect 5640 -5180 5700 -5120
rect 5740 -5180 5800 -5120
rect 5640 -5280 5700 -5220
rect 5740 -5280 5800 -5220
<< metal3 >>
rect 4000 1660 4400 1700
rect 4000 1540 4020 1660
rect 4140 1540 4260 1660
rect 4380 1540 4400 1660
rect 4000 1500 4400 1540
rect 4000 880 4200 1500
rect 4000 820 4020 880
rect 4080 820 4120 880
rect 4180 820 4200 880
rect 4000 780 4200 820
rect 4000 720 4020 780
rect 4080 720 4120 780
rect 4180 720 4200 780
rect 4000 700 4200 720
rect 1500 280 1600 300
rect 1500 220 1520 280
rect 1580 220 1600 280
rect 1500 -400 1600 220
rect 1500 -460 1520 -400
rect 1580 -460 1600 -400
rect 1500 -520 1600 -460
rect 1500 -580 1520 -520
rect 1580 -580 1600 -520
rect 1500 -1600 1600 -580
rect 1900 280 2000 300
rect 1900 220 1920 280
rect 1980 220 2000 280
rect 1900 -1300 2000 220
rect 1900 -1360 1920 -1300
rect 1980 -1360 2000 -1300
rect 1900 -1420 2000 -1360
rect 1900 -1480 1920 -1420
rect 1980 -1480 2000 -1420
rect 1900 -1600 2000 -1480
rect 2900 280 3000 300
rect 2900 220 2920 280
rect 2980 220 3000 280
rect 2900 -1300 3000 220
rect 2900 -1360 2920 -1300
rect 2980 -1360 3000 -1300
rect 2900 -1420 3000 -1360
rect 2900 -1480 2920 -1420
rect 2980 -1480 3000 -1420
rect 2900 -1600 3000 -1480
rect 3300 280 3400 300
rect 3300 220 3320 280
rect 3380 220 3400 280
rect 3300 -400 3400 220
rect 3300 -460 3320 -400
rect 3380 -460 3400 -400
rect 3300 -520 3400 -460
rect 3300 -580 3320 -520
rect 3380 -580 3400 -520
rect 3300 -1600 3400 -580
rect 5620 -5120 5820 -5100
rect 5620 -5180 5640 -5120
rect 5700 -5180 5740 -5120
rect 5800 -5180 5820 -5120
rect 5620 -5220 5820 -5180
rect 5620 -5280 5640 -5220
rect 5700 -5280 5740 -5220
rect 5800 -5280 5820 -5220
rect 5620 -5500 5820 -5280
rect 5520 -5540 5920 -5500
rect 5520 -5660 5560 -5540
rect 5680 -5660 5760 -5540
rect 5880 -5660 5920 -5540
rect 5520 -5700 5920 -5660
<< via3 >>
rect 4020 1540 4140 1660
rect 4260 1540 4380 1660
rect 5560 -5660 5680 -5540
rect 5760 -5660 5880 -5540
<< metal4 >>
rect 4000 1660 9700 1700
rect 4000 1540 4020 1660
rect 4140 1540 4260 1660
rect 4380 1540 9700 1660
rect 4000 1500 9700 1540
rect 6000 -5400 6200 1500
rect 7800 -5500 8000 1300
rect 9500 -5400 9700 1500
rect 11400 -5500 11600 1300
rect 4000 -5540 11600 -5500
rect 4000 -5660 5560 -5540
rect 5680 -5660 5760 -5540
rect 5880 -5660 11600 -5540
rect 4000 -5700 11600 -5660
use sky130_fd_pr__cap_mim_m3_1_HGK9NV  sky130_fd_pr__cap_mim_m3_1_HGK9NV_0
timestamp 1771414049
transform -1 0 9492 0 -1 -2080
box -3492 -3320 3492 3320
use sky130_fd_pr__nfet_01v8_73TUV6  sky130_fd_pr__nfet_01v8_73TUV6_0
timestamp 1771462974
transform 1 0 2088 0 1 -458
box -88 -182 88 182
use sky130_fd_pr__nfet_01v8_73TUV6  sky130_fd_pr__nfet_01v8_73TUV6_1
timestamp 1771462974
transform 1 0 2788 0 1 -458
box -88 -182 88 182
use sky130_fd_pr__nfet_01v8_73TUV6  sky130_fd_pr__nfet_01v8_73TUV6_2
timestamp 1771462974
transform 1 0 3488 0 1 -1378
box -88 -182 88 182
use sky130_fd_pr__nfet_01v8_73TUV6  sky130_fd_pr__nfet_01v8_73TUV6_3
timestamp 1771462974
transform 1 0 1388 0 1 -1378
box -88 -182 88 182
use sky130_fd_pr__nfet_01v8_K99WZJ  sky130_fd_pr__nfet_01v8_K99WZJ_0
timestamp 1771414049
transform 1 0 -1117 0 1 -603
box -183 -397 183 397
use sky130_fd_pr__nfet_01v8_PWHT78  sky130_fd_pr__nfet_01v8_PWHT78_0
timestamp 1771462974
transform 1 0 3488 0 1 -518
box -88 -182 88 182
use sky130_fd_pr__nfet_01v8_PWHT78  sky130_fd_pr__nfet_01v8_PWHT78_1
timestamp 1771462974
transform 1 0 2788 0 1 -1418
box -88 -182 88 182
use sky130_fd_pr__nfet_01v8_PWHT78  sky130_fd_pr__nfet_01v8_PWHT78_2
timestamp 1771462974
transform 1 0 2088 0 1 -1418
box -88 -182 88 182
use sky130_fd_pr__pfet_01v8_BQW8Y7  sky130_fd_pr__pfet_01v8_BQW8Y7_0
timestamp 1771462974
transform 1 0 4981 0 1 -2022
box -681 -3178 681 3144
use sky130_fd_pr__pfet_01v8_E2QEAN  sky130_fd_pr__pfet_01v8_E2QEAN_0
timestamp 1771413069
transform 1 0 -1519 0 1 734
box -681 -334 681 368
use sky130_fd_pr__res_high_po_1p41_Z9HR6K  sky130_fd_pr__res_high_po_1p41_Z9HR6K_0
timestamp 1771413069
transform 0 1 -1460 -1 0 -2019
box -141 -740 141 740
use sky130_fd_pr__res_high_po_1p41_Z9HR6K  sky130_fd_pr__res_high_po_1p41_Z9HR6K_1
timestamp 1771413069
transform 0 1 -1460 -1 0 -2359
box -141 -740 141 740
use sky130_fd_pr__res_high_po_1p41_Z9HR6K  sky130_fd_pr__res_high_po_1p41_Z9HR6K_2
timestamp 1771413069
transform 0 1 -1460 -1 0 -2699
box -141 -740 141 740
use sky130_fd_pr__res_high_po_1p41_Z9HR6K  sky130_fd_pr__res_high_po_1p41_Z9HR6K_3
timestamp 1771413069
transform 0 1 -1460 -1 0 -3039
box -141 -740 141 740
use sky130_fd_pr__nfet_01v8_PWHT78  XM2
timestamp 1771462974
transform 1 0 1388 0 1 -518
box -88 -182 88 182
use sky130_fd_pr__pfet_01v8_ES843Y  XM4
timestamp 1771413069
transform 1 0 2457 0 1 774
box -1297 -334 1297 368
use sky130_fd_pr__nfet_01v8_K99WZJ  XM5
timestamp 1771414049
transform 1 0 -517 0 1 -603
box -183 -397 183 397
use sky130_fd_pr__nfet_01v8_68987S  XM7
timestamp 1771413069
transform -1 0 3145 0 -1 -2743
box -645 -357 645 357
use sky130_fd_pr__pfet_01v8_E2QEAN  XM8
timestamp 1771413069
transform 1 0 -119 0 1 734
box -681 -334 681 368
use sky130_fd_pr__nfet_01v8_3RG5EU  XM9
timestamp 1771413069
transform 1 0 1283 0 1 -2703
box -183 -397 183 397
use sky130_fd_pr__nfet_01v8_TYFUKG  XM12
timestamp 1771413069
transform 1 0 -2027 0 1 -527
box -73 -173 73 173
use sky130_fd_pr__res_high_po_1p41_Z9HR6K  XR6
timestamp 1771413069
transform 0 1 -1460 -1 0 -1679
box -141 -740 141 740
<< labels >>
flabel metal1 40 -4580 240 -4380 0 FreeSans 256 0 0 0 VP
port 2 nsew
flabel metal1 360 -4580 560 -4380 0 FreeSans 256 0 0 0 VN
port 3 nsew
flabel metal1 -1740 1520 -1540 1720 0 FreeSans 256 0 0 0 VDD
port 0 nsew
flabel metal1 3700 -5300 3900 -5100 0 FreeSans 256 0 0 0 OUT
port 1 nsew
flabel metal1 -1540 -3800 -1340 -3600 0 FreeSans 256 0 0 0 VSS
port 4 nsew
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1771418038
<< error_p >>
rect -681 1915 681 2166
rect -681 650 681 901
rect -681 -615 681 -364
rect -681 -1880 681 -1629
rect -491 -3092 -433 -3086
rect -183 -3092 -125 -3086
rect 125 -3092 183 -3086
rect 433 -3092 491 -3086
rect -491 -3126 -479 -3092
rect -183 -3126 -171 -3092
rect 125 -3126 137 -3092
rect 433 -3126 445 -3092
rect -491 -3132 -433 -3126
rect -183 -3132 -125 -3126
rect 125 -3132 183 -3126
rect 433 -3132 491 -3126
<< nwell >>
rect -681 1915 681 3177
rect -681 650 681 1912
rect -681 -615 681 647
rect -681 -1880 681 -618
rect -681 -3145 681 -1883
<< pmos >>
rect -587 2015 -337 3115
rect -279 2015 -29 3115
rect 29 2015 279 3115
rect 337 2015 587 3115
rect -587 750 -337 1850
rect -279 750 -29 1850
rect 29 750 279 1850
rect 337 750 587 1850
rect -587 -515 -337 585
rect -279 -515 -29 585
rect 29 -515 279 585
rect 337 -515 587 585
rect -587 -1780 -337 -680
rect -279 -1780 -29 -680
rect 29 -1780 279 -680
rect 337 -1780 587 -680
rect -587 -3045 -337 -1945
rect -279 -3045 -29 -1945
rect 29 -3045 279 -1945
rect 337 -3045 587 -1945
<< pdiff >>
rect -645 2834 -587 3115
rect -645 2296 -633 2834
rect -599 2296 -587 2834
rect -645 2015 -587 2296
rect -337 2834 -279 3115
rect -337 2296 -325 2834
rect -291 2296 -279 2834
rect -337 2015 -279 2296
rect -29 2834 29 3115
rect -29 2296 -17 2834
rect 17 2296 29 2834
rect -29 2015 29 2296
rect 279 2834 337 3115
rect 279 2296 291 2834
rect 325 2296 337 2834
rect 279 2015 337 2296
rect 587 2834 645 3115
rect 587 2296 599 2834
rect 633 2296 645 2834
rect 587 2015 645 2296
rect -645 1569 -587 1850
rect -645 1031 -633 1569
rect -599 1031 -587 1569
rect -645 750 -587 1031
rect -337 1569 -279 1850
rect -337 1031 -325 1569
rect -291 1031 -279 1569
rect -337 750 -279 1031
rect -29 1569 29 1850
rect -29 1031 -17 1569
rect 17 1031 29 1569
rect -29 750 29 1031
rect 279 1569 337 1850
rect 279 1031 291 1569
rect 325 1031 337 1569
rect 279 750 337 1031
rect 587 1569 645 1850
rect 587 1031 599 1569
rect 633 1031 645 1569
rect 587 750 645 1031
rect -645 304 -587 585
rect -645 -234 -633 304
rect -599 -234 -587 304
rect -645 -515 -587 -234
rect -337 304 -279 585
rect -337 -234 -325 304
rect -291 -234 -279 304
rect -337 -515 -279 -234
rect -29 304 29 585
rect -29 -234 -17 304
rect 17 -234 29 304
rect -29 -515 29 -234
rect 279 304 337 585
rect 279 -234 291 304
rect 325 -234 337 304
rect 279 -515 337 -234
rect 587 304 645 585
rect 587 -234 599 304
rect 633 -234 645 304
rect 587 -515 645 -234
rect -645 -961 -587 -680
rect -645 -1499 -633 -961
rect -599 -1499 -587 -961
rect -645 -1780 -587 -1499
rect -337 -961 -279 -680
rect -337 -1499 -325 -961
rect -291 -1499 -279 -961
rect -337 -1780 -279 -1499
rect -29 -961 29 -680
rect -29 -1499 -17 -961
rect 17 -1499 29 -961
rect -29 -1780 29 -1499
rect 279 -961 337 -680
rect 279 -1499 291 -961
rect 325 -1499 337 -961
rect 279 -1780 337 -1499
rect 587 -961 645 -680
rect 587 -1499 599 -961
rect 633 -1499 645 -961
rect 587 -1780 645 -1499
rect -645 -2226 -587 -1945
rect -645 -2764 -633 -2226
rect -599 -2764 -587 -2226
rect -645 -3045 -587 -2764
rect -337 -2226 -279 -1945
rect -337 -2764 -325 -2226
rect -291 -2764 -279 -2226
rect -337 -3045 -279 -2764
rect -29 -2226 29 -1945
rect -29 -2764 -17 -2226
rect 17 -2764 29 -2226
rect -29 -3045 29 -2764
rect 279 -2226 337 -1945
rect 279 -2764 291 -2226
rect 325 -2764 337 -2226
rect 279 -3045 337 -2764
rect 587 -2226 645 -1945
rect 587 -2764 599 -2226
rect 633 -2764 645 -2226
rect 587 -3045 645 -2764
<< pdiffc >>
rect -633 2296 -599 2834
rect -325 2296 -291 2834
rect -17 2296 17 2834
rect 291 2296 325 2834
rect 599 2296 633 2834
rect -633 1031 -599 1569
rect -325 1031 -291 1569
rect -17 1031 17 1569
rect 291 1031 325 1569
rect 599 1031 633 1569
rect -633 -234 -599 304
rect -325 -234 -291 304
rect -17 -234 17 304
rect 291 -234 325 304
rect 599 -234 633 304
rect -633 -1499 -599 -961
rect -325 -1499 -291 -961
rect -17 -1499 17 -961
rect 291 -1499 325 -961
rect 599 -1499 633 -961
rect -633 -2764 -599 -2226
rect -325 -2764 -291 -2226
rect -17 -2764 17 -2226
rect 291 -2764 325 -2226
rect 599 -2764 633 -2226
<< poly >>
rect -587 3115 -337 3141
rect -279 3115 -29 3141
rect 29 3115 279 3141
rect 337 3115 587 3141
rect -587 1968 -337 2015
rect -587 1951 -484 1968
rect -500 1934 -484 1951
rect -440 1951 -337 1968
rect -279 1968 -29 2015
rect -279 1951 -176 1968
rect -440 1934 -424 1951
rect -500 1918 -424 1934
rect -192 1934 -176 1951
rect -132 1951 -29 1968
rect 29 1968 279 2015
rect 29 1951 132 1968
rect -132 1934 -116 1951
rect -192 1918 -116 1934
rect 116 1934 132 1951
rect 176 1951 279 1968
rect 337 1968 587 2015
rect 337 1951 440 1968
rect 176 1934 192 1951
rect 116 1918 192 1934
rect 424 1934 440 1951
rect 484 1951 587 1968
rect 484 1934 500 1951
rect 424 1918 500 1934
rect -587 1850 -337 1876
rect -279 1850 -29 1876
rect 29 1850 279 1876
rect 337 1850 587 1876
rect -587 703 -337 750
rect -587 686 -484 703
rect -500 669 -484 686
rect -440 686 -337 703
rect -279 703 -29 750
rect -279 686 -176 703
rect -440 669 -424 686
rect -500 653 -424 669
rect -192 669 -176 686
rect -132 686 -29 703
rect 29 703 279 750
rect 29 686 132 703
rect -132 669 -116 686
rect -192 653 -116 669
rect 116 669 132 686
rect 176 686 279 703
rect 337 703 587 750
rect 337 686 440 703
rect 176 669 192 686
rect 116 653 192 669
rect 424 669 440 686
rect 484 686 587 703
rect 484 669 500 686
rect 424 653 500 669
rect -587 585 -337 611
rect -279 585 -29 611
rect 29 585 279 611
rect 337 585 587 611
rect -587 -562 -337 -515
rect -587 -579 -484 -562
rect -500 -596 -484 -579
rect -440 -579 -337 -562
rect -279 -562 -29 -515
rect -279 -579 -176 -562
rect -440 -596 -424 -579
rect -500 -612 -424 -596
rect -192 -596 -176 -579
rect -132 -579 -29 -562
rect 29 -562 279 -515
rect 29 -579 132 -562
rect -132 -596 -116 -579
rect -192 -612 -116 -596
rect 116 -596 132 -579
rect 176 -579 279 -562
rect 337 -562 587 -515
rect 337 -579 440 -562
rect 176 -596 192 -579
rect 116 -612 192 -596
rect 424 -596 440 -579
rect 484 -579 587 -562
rect 484 -596 500 -579
rect 424 -612 500 -596
rect -587 -680 -337 -654
rect -279 -680 -29 -654
rect 29 -680 279 -654
rect 337 -680 587 -654
rect -587 -1827 -337 -1780
rect -587 -1844 -484 -1827
rect -500 -1861 -484 -1844
rect -440 -1844 -337 -1827
rect -279 -1827 -29 -1780
rect -279 -1844 -176 -1827
rect -440 -1861 -424 -1844
rect -500 -1877 -424 -1861
rect -192 -1861 -176 -1844
rect -132 -1844 -29 -1827
rect 29 -1827 279 -1780
rect 29 -1844 132 -1827
rect -132 -1861 -116 -1844
rect -192 -1877 -116 -1861
rect 116 -1861 132 -1844
rect 176 -1844 279 -1827
rect 337 -1827 587 -1780
rect 337 -1844 440 -1827
rect 176 -1861 192 -1844
rect 116 -1877 192 -1861
rect 424 -1861 440 -1844
rect 484 -1844 587 -1827
rect 484 -1861 500 -1844
rect 424 -1877 500 -1861
rect -587 -1945 -337 -1919
rect -279 -1945 -29 -1919
rect 29 -1945 279 -1919
rect 337 -1945 587 -1919
rect -587 -3092 -337 -3045
rect -587 -3109 -484 -3092
rect -500 -3126 -484 -3109
rect -440 -3109 -337 -3092
rect -279 -3092 -29 -3045
rect -279 -3109 -176 -3092
rect -440 -3126 -424 -3109
rect -500 -3142 -424 -3126
rect -192 -3126 -176 -3109
rect -132 -3109 -29 -3092
rect 29 -3092 279 -3045
rect 29 -3109 132 -3092
rect -132 -3126 -116 -3109
rect -192 -3142 -116 -3126
rect 116 -3126 132 -3109
rect 176 -3109 279 -3092
rect 337 -3092 587 -3045
rect 337 -3109 440 -3092
rect 176 -3126 192 -3109
rect 116 -3142 192 -3126
rect 424 -3126 440 -3109
rect 484 -3109 587 -3092
rect 484 -3126 500 -3109
rect 424 -3142 500 -3126
<< polycont >>
rect -484 1934 -440 1968
rect -176 1934 -132 1968
rect 132 1934 176 1968
rect 440 1934 484 1968
rect -484 669 -440 703
rect -176 669 -132 703
rect 132 669 176 703
rect 440 669 484 703
rect -484 -596 -440 -562
rect -176 -596 -132 -562
rect 132 -596 176 -562
rect 440 -596 484 -562
rect -484 -1861 -440 -1827
rect -176 -1861 -132 -1827
rect 132 -1861 176 -1827
rect 440 -1861 484 -1827
rect -484 -3126 -440 -3092
rect -176 -3126 -132 -3092
rect 132 -3126 176 -3092
rect 440 -3126 484 -3092
<< locali >>
rect -633 2834 -599 2850
rect -633 2280 -599 2296
rect -325 2834 -291 2850
rect -325 2280 -291 2296
rect -17 2834 17 2850
rect -17 2280 17 2296
rect 291 2834 325 2850
rect 291 2280 325 2296
rect 599 2834 633 2850
rect 599 2280 633 2296
rect -500 1934 -484 1968
rect -440 1934 -424 1968
rect -192 1934 -176 1968
rect -132 1934 -116 1968
rect 116 1934 132 1968
rect 176 1934 192 1968
rect 424 1934 440 1968
rect 484 1934 500 1968
rect -633 1569 -599 1585
rect -633 1015 -599 1031
rect -325 1569 -291 1585
rect -325 1015 -291 1031
rect -17 1569 17 1585
rect -17 1015 17 1031
rect 291 1569 325 1585
rect 291 1015 325 1031
rect 599 1569 633 1585
rect 599 1015 633 1031
rect -500 669 -484 703
rect -440 669 -424 703
rect -192 669 -176 703
rect -132 669 -116 703
rect 116 669 132 703
rect 176 669 192 703
rect 424 669 440 703
rect 484 669 500 703
rect -633 304 -599 320
rect -633 -250 -599 -234
rect -325 304 -291 320
rect -325 -250 -291 -234
rect -17 304 17 320
rect -17 -250 17 -234
rect 291 304 325 320
rect 291 -250 325 -234
rect 599 304 633 320
rect 599 -250 633 -234
rect -500 -596 -484 -562
rect -440 -596 -424 -562
rect -192 -596 -176 -562
rect -132 -596 -116 -562
rect 116 -596 132 -562
rect 176 -596 192 -562
rect 424 -596 440 -562
rect 484 -596 500 -562
rect -633 -961 -599 -945
rect -633 -1515 -599 -1499
rect -325 -961 -291 -945
rect -325 -1515 -291 -1499
rect -17 -961 17 -945
rect -17 -1515 17 -1499
rect 291 -961 325 -945
rect 291 -1515 325 -1499
rect 599 -961 633 -945
rect 599 -1515 633 -1499
rect -500 -1861 -484 -1827
rect -440 -1861 -424 -1827
rect -192 -1861 -176 -1827
rect -132 -1861 -116 -1827
rect 116 -1861 132 -1827
rect 176 -1861 192 -1827
rect 424 -1861 440 -1827
rect 484 -1861 500 -1827
rect -633 -2226 -599 -2210
rect -633 -2780 -599 -2764
rect -325 -2226 -291 -2210
rect -325 -2780 -291 -2764
rect -17 -2226 17 -2210
rect -17 -2780 17 -2764
rect 291 -2226 325 -2210
rect 291 -2780 325 -2764
rect 599 -2226 633 -2210
rect 599 -2780 633 -2764
rect -500 -3126 -484 -3092
rect -440 -3126 -424 -3092
rect -192 -3126 -176 -3092
rect -132 -3126 -116 -3092
rect 116 -3126 132 -3092
rect 176 -3126 192 -3092
rect 424 -3126 440 -3092
rect 484 -3126 500 -3092
<< viali >>
rect -633 2296 -599 2834
rect -325 2296 -291 2834
rect -17 2296 17 2834
rect 291 2296 325 2834
rect 599 2296 633 2834
rect -479 1934 -445 1968
rect -171 1934 -137 1968
rect 137 1934 171 1968
rect 445 1934 479 1968
rect -633 1031 -599 1569
rect -325 1031 -291 1569
rect -17 1031 17 1569
rect 291 1031 325 1569
rect 599 1031 633 1569
rect -479 669 -445 703
rect -171 669 -137 703
rect 137 669 171 703
rect 445 669 479 703
rect -633 -234 -599 304
rect -325 -234 -291 304
rect -17 -234 17 304
rect 291 -234 325 304
rect 599 -234 633 304
rect -479 -596 -445 -562
rect -171 -596 -137 -562
rect 137 -596 171 -562
rect 445 -596 479 -562
rect -633 -1499 -599 -961
rect -325 -1499 -291 -961
rect -17 -1499 17 -961
rect 291 -1499 325 -961
rect 599 -1499 633 -961
rect -479 -1861 -445 -1827
rect -171 -1861 -137 -1827
rect 137 -1861 171 -1827
rect 445 -1861 479 -1827
rect -633 -2764 -599 -2226
rect -325 -2764 -291 -2226
rect -17 -2764 17 -2226
rect 291 -2764 325 -2226
rect 599 -2764 633 -2226
rect -479 -3126 -445 -3092
rect -171 -3126 -137 -3092
rect 137 -3126 171 -3092
rect 445 -3126 479 -3092
<< metal1 >>
rect -639 2834 -593 2846
rect -639 2296 -633 2834
rect -599 2296 -593 2834
rect -639 2284 -593 2296
rect -331 2834 -285 2846
rect -331 2296 -325 2834
rect -291 2296 -285 2834
rect -331 2284 -285 2296
rect -23 2834 23 2846
rect -23 2296 -17 2834
rect 17 2296 23 2834
rect -23 2284 23 2296
rect 285 2834 331 2846
rect 285 2296 291 2834
rect 325 2296 331 2834
rect 285 2284 331 2296
rect 593 2834 639 2846
rect 593 2296 599 2834
rect 633 2296 639 2834
rect 593 2284 639 2296
rect -491 1968 -433 1974
rect -491 1934 -479 1968
rect -445 1934 -433 1968
rect -491 1928 -433 1934
rect -183 1968 -125 1974
rect -183 1934 -171 1968
rect -137 1934 -125 1968
rect -183 1928 -125 1934
rect 125 1968 183 1974
rect 125 1934 137 1968
rect 171 1934 183 1968
rect 125 1928 183 1934
rect 433 1968 491 1974
rect 433 1934 445 1968
rect 479 1934 491 1968
rect 433 1928 491 1934
rect -639 1569 -593 1581
rect -639 1031 -633 1569
rect -599 1031 -593 1569
rect -639 1019 -593 1031
rect -331 1569 -285 1581
rect -331 1031 -325 1569
rect -291 1031 -285 1569
rect -331 1019 -285 1031
rect -23 1569 23 1581
rect -23 1031 -17 1569
rect 17 1031 23 1569
rect -23 1019 23 1031
rect 285 1569 331 1581
rect 285 1031 291 1569
rect 325 1031 331 1569
rect 285 1019 331 1031
rect 593 1569 639 1581
rect 593 1031 599 1569
rect 633 1031 639 1569
rect 593 1019 639 1031
rect -491 703 -433 709
rect -491 669 -479 703
rect -445 669 -433 703
rect -491 663 -433 669
rect -183 703 -125 709
rect -183 669 -171 703
rect -137 669 -125 703
rect -183 663 -125 669
rect 125 703 183 709
rect 125 669 137 703
rect 171 669 183 703
rect 125 663 183 669
rect 433 703 491 709
rect 433 669 445 703
rect 479 669 491 703
rect 433 663 491 669
rect -639 304 -593 316
rect -639 -234 -633 304
rect -599 -234 -593 304
rect -639 -246 -593 -234
rect -331 304 -285 316
rect -331 -234 -325 304
rect -291 -234 -285 304
rect -331 -246 -285 -234
rect -23 304 23 316
rect -23 -234 -17 304
rect 17 -234 23 304
rect -23 -246 23 -234
rect 285 304 331 316
rect 285 -234 291 304
rect 325 -234 331 304
rect 285 -246 331 -234
rect 593 304 639 316
rect 593 -234 599 304
rect 633 -234 639 304
rect 593 -246 639 -234
rect -491 -562 -433 -556
rect -491 -596 -479 -562
rect -445 -596 -433 -562
rect -491 -602 -433 -596
rect -183 -562 -125 -556
rect -183 -596 -171 -562
rect -137 -596 -125 -562
rect -183 -602 -125 -596
rect 125 -562 183 -556
rect 125 -596 137 -562
rect 171 -596 183 -562
rect 125 -602 183 -596
rect 433 -562 491 -556
rect 433 -596 445 -562
rect 479 -596 491 -562
rect 433 -602 491 -596
rect -639 -961 -593 -949
rect -639 -1499 -633 -961
rect -599 -1499 -593 -961
rect -639 -1511 -593 -1499
rect -331 -961 -285 -949
rect -331 -1499 -325 -961
rect -291 -1499 -285 -961
rect -331 -1511 -285 -1499
rect -23 -961 23 -949
rect -23 -1499 -17 -961
rect 17 -1499 23 -961
rect -23 -1511 23 -1499
rect 285 -961 331 -949
rect 285 -1499 291 -961
rect 325 -1499 331 -961
rect 285 -1511 331 -1499
rect 593 -961 639 -949
rect 593 -1499 599 -961
rect 633 -1499 639 -961
rect 593 -1511 639 -1499
rect -491 -1827 -433 -1821
rect -491 -1861 -479 -1827
rect -445 -1861 -433 -1827
rect -491 -1867 -433 -1861
rect -183 -1827 -125 -1821
rect -183 -1861 -171 -1827
rect -137 -1861 -125 -1827
rect -183 -1867 -125 -1861
rect 125 -1827 183 -1821
rect 125 -1861 137 -1827
rect 171 -1861 183 -1827
rect 125 -1867 183 -1861
rect 433 -1827 491 -1821
rect 433 -1861 445 -1827
rect 479 -1861 491 -1827
rect 433 -1867 491 -1861
rect -639 -2226 -593 -2214
rect -639 -2764 -633 -2226
rect -599 -2764 -593 -2226
rect -639 -2776 -593 -2764
rect -331 -2226 -285 -2214
rect -331 -2764 -325 -2226
rect -291 -2764 -285 -2226
rect -331 -2776 -285 -2764
rect -23 -2226 23 -2214
rect -23 -2764 -17 -2226
rect 17 -2764 23 -2226
rect -23 -2776 23 -2764
rect 285 -2226 331 -2214
rect 285 -2764 291 -2226
rect 325 -2764 331 -2226
rect 285 -2776 331 -2764
rect 593 -2226 639 -2214
rect 593 -2764 599 -2226
rect 633 -2764 639 -2226
rect 593 -2776 639 -2764
rect -491 -3092 -433 -3086
rect -491 -3126 -479 -3092
rect -445 -3126 -433 -3092
rect -491 -3132 -433 -3126
rect -183 -3092 -125 -3086
rect -183 -3126 -171 -3092
rect -137 -3126 -125 -3092
rect -183 -3132 -125 -3126
rect 125 -3092 183 -3086
rect 125 -3126 137 -3092
rect 171 -3126 183 -3092
rect 125 -3132 183 -3126
rect 433 -3092 491 -3086
rect 433 -3126 445 -3092
rect 479 -3126 491 -3092
rect 433 -3132 491 -3126
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 5.5 l 1.25 m 5 nf 4 diffcov 50 polycov 20 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 class mosfet compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 50 viadrn 50 viagate 10 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1770979109
<< nwell >>
rect -2283 -944 2283 944
<< pmos >>
rect -2087 -725 -1087 725
rect -1029 -725 -29 725
rect 29 -725 1029 725
rect 1087 -725 2087 725
<< pdiff >>
rect -2145 713 -2087 725
rect -2145 -713 -2133 713
rect -2099 -713 -2087 713
rect -2145 -725 -2087 -713
rect -1087 713 -1029 725
rect -1087 -713 -1075 713
rect -1041 -713 -1029 713
rect -1087 -725 -1029 -713
rect -29 713 29 725
rect -29 -713 -17 713
rect 17 -713 29 713
rect -29 -725 29 -713
rect 1029 713 1087 725
rect 1029 -713 1041 713
rect 1075 -713 1087 713
rect 1029 -725 1087 -713
rect 2087 713 2145 725
rect 2087 -713 2099 713
rect 2133 -713 2145 713
rect 2087 -725 2145 -713
<< pdiffc >>
rect -2133 -713 -2099 713
rect -1075 -713 -1041 713
rect -17 -713 17 713
rect 1041 -713 1075 713
rect 2099 -713 2133 713
<< nsubdiff >>
rect -2247 874 -2151 908
rect 2151 874 2247 908
rect -2247 812 -2213 874
rect 2213 812 2247 874
rect -2247 -874 -2213 -812
rect 2213 -874 2247 -812
rect -2247 -908 -2151 -874
rect 2151 -908 2247 -874
<< nsubdiffcont >>
rect -2151 874 2151 908
rect -2247 -812 -2213 812
rect 2213 -812 2247 812
rect -2151 -908 2151 -874
<< poly >>
rect -2087 806 -1087 822
rect -2087 772 -2071 806
rect -1103 772 -1087 806
rect -2087 725 -1087 772
rect -1029 806 -29 822
rect -1029 772 -1013 806
rect -45 772 -29 806
rect -1029 725 -29 772
rect 29 806 1029 822
rect 29 772 45 806
rect 1013 772 1029 806
rect 29 725 1029 772
rect 1087 806 2087 822
rect 1087 772 1103 806
rect 2071 772 2087 806
rect 1087 725 2087 772
rect -2087 -772 -1087 -725
rect -2087 -806 -2071 -772
rect -1103 -806 -1087 -772
rect -2087 -822 -1087 -806
rect -1029 -772 -29 -725
rect -1029 -806 -1013 -772
rect -45 -806 -29 -772
rect -1029 -822 -29 -806
rect 29 -772 1029 -725
rect 29 -806 45 -772
rect 1013 -806 1029 -772
rect 29 -822 1029 -806
rect 1087 -772 2087 -725
rect 1087 -806 1103 -772
rect 2071 -806 2087 -772
rect 1087 -822 2087 -806
<< polycont >>
rect -2071 772 -1103 806
rect -1013 772 -45 806
rect 45 772 1013 806
rect 1103 772 2071 806
rect -2071 -806 -1103 -772
rect -1013 -806 -45 -772
rect 45 -806 1013 -772
rect 1103 -806 2071 -772
<< locali >>
rect -2247 874 -2151 908
rect 2151 874 2247 908
rect -2247 812 -2213 874
rect 2213 812 2247 874
rect -2087 772 -2071 806
rect -1103 772 -1087 806
rect -1029 772 -1013 806
rect -45 772 -29 806
rect 29 772 45 806
rect 1013 772 1029 806
rect 1087 772 1103 806
rect 2071 772 2087 806
rect -2133 713 -2099 729
rect -2133 -729 -2099 -713
rect -1075 713 -1041 729
rect -1075 -729 -1041 -713
rect -17 713 17 729
rect -17 -729 17 -713
rect 1041 713 1075 729
rect 1041 -729 1075 -713
rect 2099 713 2133 729
rect 2099 -729 2133 -713
rect -2087 -806 -2071 -772
rect -1103 -806 -1087 -772
rect -1029 -806 -1013 -772
rect -45 -806 -29 -772
rect 29 -806 45 -772
rect 1013 -806 1029 -772
rect 1087 -806 1103 -772
rect 2071 -806 2087 -772
rect -2247 -874 -2213 -812
rect 2213 -874 2247 -812
rect -2247 -908 -2151 -874
rect 2151 -908 2247 -874
<< viali >>
rect -2071 772 -1103 806
rect -1013 772 -45 806
rect 45 772 1013 806
rect 1103 772 2071 806
rect -2133 -713 -2099 713
rect -1075 -713 -1041 713
rect -17 -713 17 713
rect 1041 -713 1075 713
rect 2099 -713 2133 713
rect -2071 -806 -1103 -772
rect -1013 -806 -45 -772
rect 45 -806 1013 -772
rect 1103 -806 2071 -772
<< metal1 >>
rect -2083 806 -1091 812
rect -2083 772 -2071 806
rect -1103 772 -1091 806
rect -2083 766 -1091 772
rect -1025 806 -33 812
rect -1025 772 -1013 806
rect -45 772 -33 806
rect -1025 766 -33 772
rect 33 806 1025 812
rect 33 772 45 806
rect 1013 772 1025 806
rect 33 766 1025 772
rect 1091 806 2083 812
rect 1091 772 1103 806
rect 2071 772 2083 806
rect 1091 766 2083 772
rect -2139 713 -2093 725
rect -2139 -713 -2133 713
rect -2099 -713 -2093 713
rect -2139 -725 -2093 -713
rect -1081 713 -1035 725
rect -1081 -713 -1075 713
rect -1041 -713 -1035 713
rect -1081 -725 -1035 -713
rect -23 713 23 725
rect -23 -713 -17 713
rect 17 -713 23 713
rect -23 -725 23 -713
rect 1035 713 1081 725
rect 1035 -713 1041 713
rect 1075 -713 1081 713
rect 1035 -725 1081 -713
rect 2093 713 2139 725
rect 2093 -713 2099 713
rect 2133 -713 2139 713
rect 2093 -725 2139 -713
rect -2083 -772 -1091 -766
rect -2083 -806 -2071 -772
rect -1103 -806 -1091 -772
rect -2083 -812 -1091 -806
rect -1025 -772 -33 -766
rect -1025 -806 -1013 -772
rect -45 -806 -33 -772
rect -1025 -812 -33 -806
rect 33 -772 1025 -766
rect 33 -806 45 -772
rect 1013 -806 1025 -772
rect 33 -812 1025 -806
rect 1091 -772 2083 -766
rect 1091 -806 1103 -772
rect 2071 -806 2083 -772
rect 1091 -812 2083 -806
<< properties >>
string FIXED_BBOX -2230 -891 2230 891
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 7.25 l 5.0 m 1 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 class mosfet compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1771413069
<< nwell >>
rect -1297 -370 1297 370
<< pmos >>
rect -1203 -270 -953 270
rect -895 -270 -645 270
rect -587 -270 -337 270
rect -279 -270 -29 270
rect 29 -270 279 270
rect 337 -270 587 270
rect 645 -270 895 270
rect 953 -270 1203 270
<< pdiff >>
rect -1261 258 -1203 270
rect -1261 -258 -1249 258
rect -1215 -258 -1203 258
rect -1261 -270 -1203 -258
rect -953 258 -895 270
rect -953 -258 -941 258
rect -907 -258 -895 258
rect -953 -270 -895 -258
rect -645 258 -587 270
rect -645 -258 -633 258
rect -599 -258 -587 258
rect -645 -270 -587 -258
rect -337 258 -279 270
rect -337 -258 -325 258
rect -291 -258 -279 258
rect -337 -270 -279 -258
rect -29 258 29 270
rect -29 -258 -17 258
rect 17 -258 29 258
rect -29 -270 29 -258
rect 279 258 337 270
rect 279 -258 291 258
rect 325 -258 337 258
rect 279 -270 337 -258
rect 587 258 645 270
rect 587 -258 599 258
rect 633 -258 645 258
rect 587 -270 645 -258
rect 895 258 953 270
rect 895 -258 907 258
rect 941 -258 953 258
rect 895 -270 953 -258
rect 1203 258 1261 270
rect 1203 -258 1215 258
rect 1249 -258 1261 258
rect 1203 -270 1261 -258
<< pdiffc >>
rect -1249 -258 -1215 258
rect -941 -258 -907 258
rect -633 -258 -599 258
rect -325 -258 -291 258
rect -17 -258 17 258
rect 291 -258 325 258
rect 599 -258 633 258
rect 907 -258 941 258
rect 1215 -258 1249 258
<< poly >>
rect -1203 351 -953 367
rect -1203 317 -1187 351
rect -969 317 -953 351
rect -1203 270 -953 317
rect -895 351 -645 367
rect -895 317 -879 351
rect -661 317 -645 351
rect -895 270 -645 317
rect -587 351 -337 367
rect -587 317 -571 351
rect -353 317 -337 351
rect -587 270 -337 317
rect -279 351 -29 367
rect -279 317 -263 351
rect -45 317 -29 351
rect -279 270 -29 317
rect 29 351 279 367
rect 29 317 45 351
rect 263 317 279 351
rect 29 270 279 317
rect 337 351 587 367
rect 337 317 353 351
rect 571 317 587 351
rect 337 270 587 317
rect 645 351 895 367
rect 645 317 661 351
rect 879 317 895 351
rect 645 270 895 317
rect 953 351 1203 367
rect 953 317 969 351
rect 1187 317 1203 351
rect 953 270 1203 317
rect -1203 -317 -953 -270
rect -1203 -351 -1187 -317
rect -969 -351 -953 -317
rect -1203 -367 -953 -351
rect -895 -317 -645 -270
rect -895 -351 -879 -317
rect -661 -351 -645 -317
rect -895 -367 -645 -351
rect -587 -317 -337 -270
rect -587 -351 -571 -317
rect -353 -351 -337 -317
rect -587 -367 -337 -351
rect -279 -317 -29 -270
rect -279 -351 -263 -317
rect -45 -351 -29 -317
rect -279 -367 -29 -351
rect 29 -317 279 -270
rect 29 -351 45 -317
rect 263 -351 279 -317
rect 29 -367 279 -351
rect 337 -317 587 -270
rect 337 -351 353 -317
rect 571 -351 587 -317
rect 337 -367 587 -351
rect 645 -317 895 -270
rect 645 -351 661 -317
rect 879 -351 895 -317
rect 645 -367 895 -351
rect 953 -317 1203 -270
rect 953 -351 969 -317
rect 1187 -351 1203 -317
rect 953 -367 1203 -351
<< polycont >>
rect -1187 317 -969 351
rect -879 317 -661 351
rect -571 317 -353 351
rect -263 317 -45 351
rect 45 317 263 351
rect 353 317 571 351
rect 661 317 879 351
rect 969 317 1187 351
rect -1187 -351 -969 -317
rect -879 -351 -661 -317
rect -571 -351 -353 -317
rect -263 -351 -45 -317
rect 45 -351 263 -317
rect 353 -351 571 -317
rect 661 -351 879 -317
rect 969 -351 1187 -317
<< locali >>
rect -1203 317 -1187 351
rect -969 317 -953 351
rect -895 317 -879 351
rect -661 317 -645 351
rect -587 317 -571 351
rect -353 317 -337 351
rect -279 317 -263 351
rect -45 317 -29 351
rect 29 317 45 351
rect 263 317 279 351
rect 337 317 353 351
rect 571 317 587 351
rect 645 317 661 351
rect 879 317 895 351
rect 953 317 969 351
rect 1187 317 1203 351
rect -1249 258 -1215 274
rect -1249 -274 -1215 -258
rect -941 258 -907 274
rect -941 -274 -907 -258
rect -633 258 -599 274
rect -633 -274 -599 -258
rect -325 258 -291 274
rect -325 -274 -291 -258
rect -17 258 17 274
rect -17 -274 17 -258
rect 291 258 325 274
rect 291 -274 325 -258
rect 599 258 633 274
rect 599 -274 633 -258
rect 907 258 941 274
rect 907 -274 941 -258
rect 1215 258 1249 274
rect 1215 -274 1249 -258
rect -1203 -351 -1187 -317
rect -969 -351 -953 -317
rect -895 -351 -879 -317
rect -661 -351 -645 -317
rect -587 -351 -571 -317
rect -353 -351 -337 -317
rect -279 -351 -263 -317
rect -45 -351 -29 -317
rect 29 -351 45 -317
rect 263 -351 279 -317
rect 337 -351 353 -317
rect 571 -351 587 -317
rect 645 -351 661 -317
rect 879 -351 895 -317
rect 953 -351 969 -317
rect 1187 -351 1203 -317
<< viali >>
rect -1187 317 -969 351
rect -879 317 -661 351
rect -571 317 -353 351
rect -263 317 -45 351
rect 45 317 263 351
rect 353 317 571 351
rect 661 317 879 351
rect 969 317 1187 351
rect -1249 -258 -1215 258
rect -941 -258 -907 258
rect -633 -258 -599 258
rect -325 -258 -291 258
rect -17 -258 17 258
rect 291 -258 325 258
rect 599 -258 633 258
rect 907 -258 941 258
rect 1215 -258 1249 258
rect -1187 -351 -969 -317
rect -879 -351 -661 -317
rect -571 -351 -353 -317
rect -263 -351 -45 -317
rect 45 -351 263 -317
rect 353 -351 571 -317
rect 661 -351 879 -317
rect 969 -351 1187 -317
<< metal1 >>
rect -1199 351 -957 357
rect -1199 317 -1187 351
rect -969 317 -957 351
rect -1199 311 -957 317
rect -891 351 -649 357
rect -891 317 -879 351
rect -661 317 -649 351
rect -891 311 -649 317
rect -583 351 -341 357
rect -583 317 -571 351
rect -353 317 -341 351
rect -583 311 -341 317
rect -275 351 -33 357
rect -275 317 -263 351
rect -45 317 -33 351
rect -275 311 -33 317
rect 33 351 275 357
rect 33 317 45 351
rect 263 317 275 351
rect 33 311 275 317
rect 341 351 583 357
rect 341 317 353 351
rect 571 317 583 351
rect 341 311 583 317
rect 649 351 891 357
rect 649 317 661 351
rect 879 317 891 351
rect 649 311 891 317
rect 957 351 1199 357
rect 957 317 969 351
rect 1187 317 1199 351
rect 957 311 1199 317
rect -1255 258 -1209 270
rect -1255 -258 -1249 258
rect -1215 -258 -1209 258
rect -1255 -270 -1209 -258
rect -947 258 -901 270
rect -947 -258 -941 258
rect -907 -258 -901 258
rect -947 -270 -901 -258
rect -639 258 -593 270
rect -639 -258 -633 258
rect -599 -258 -593 258
rect -639 -270 -593 -258
rect -331 258 -285 270
rect -331 -258 -325 258
rect -291 -258 -285 258
rect -331 -270 -285 -258
rect -23 258 23 270
rect -23 -258 -17 258
rect 17 -258 23 258
rect -23 -270 23 -258
rect 285 258 331 270
rect 285 -258 291 258
rect 325 -258 331 258
rect 285 -270 331 -258
rect 593 258 639 270
rect 593 -258 599 258
rect 633 -258 639 258
rect 593 -270 639 -258
rect 901 258 947 270
rect 901 -258 907 258
rect 941 -258 947 258
rect 901 -270 947 -258
rect 1209 258 1255 270
rect 1209 -258 1215 258
rect 1249 -258 1255 258
rect 1209 -270 1255 -258
rect -1199 -317 -957 -311
rect -1199 -351 -1187 -317
rect -969 -351 -957 -317
rect -1199 -357 -957 -351
rect -891 -317 -649 -311
rect -891 -351 -879 -317
rect -661 -351 -649 -317
rect -891 -357 -649 -351
rect -583 -317 -341 -311
rect -583 -351 -571 -317
rect -353 -351 -341 -317
rect -583 -357 -341 -351
rect -275 -317 -33 -311
rect -275 -351 -263 -317
rect -45 -351 -33 -317
rect -275 -357 -33 -351
rect 33 -317 275 -311
rect 33 -351 45 -317
rect 263 -351 275 -317
rect 33 -357 275 -351
rect 341 -317 583 -311
rect 341 -351 353 -317
rect 571 -351 583 -317
rect 341 -357 583 -351
rect 649 -317 891 -311
rect 649 -351 661 -317
rect 879 -351 891 -317
rect 649 -357 891 -351
rect 957 -317 1199 -311
rect 957 -351 969 -317
rect 1187 -351 1199 -317
rect 957 -357 1199 -351
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 2.7 l 1.25 m 1 nf 8 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 class mosfet compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1771083444
<< nwell >>
rect -1660 2040 9860 4040
rect -1660 -2560 1460 2040
rect 6740 -2560 9860 2040
rect -1660 -4660 9860 -2560
<< pwell >>
rect 1500 -840 6700 2000
rect 1500 -900 2360 -840
rect 2380 -900 5880 -840
rect 5900 -900 6700 -840
rect 1500 -2350 6700 -900
rect 1500 -2360 2280 -2350
rect 5980 -2360 6700 -2350
rect 1500 -2400 6700 -2360
rect 1500 -2510 6700 -2410
<< psubdiff >>
rect 1500 1980 6700 2000
rect 1500 1920 1620 1980
rect 6580 1920 6700 1980
rect 1500 1900 6700 1920
rect 1500 1880 1600 1900
rect 1500 -2380 1520 1880
rect 1580 -2380 1600 1880
rect 6600 1880 6700 1900
rect 1700 1780 6500 1800
rect 1700 1720 1820 1780
rect 6380 1720 6500 1780
rect 1700 1700 6500 1720
rect 1700 1680 1800 1700
rect 1700 320 1720 1680
rect 1780 320 1800 1680
rect 1700 300 1800 320
rect 6400 1680 6500 1700
rect 6400 320 6420 1680
rect 6480 320 6500 1680
rect 6400 300 6500 320
rect 1700 280 6500 300
rect 1700 220 1820 280
rect 3040 220 5160 280
rect 6380 220 6500 280
rect 1700 200 6500 220
rect 1700 80 2800 100
rect 1700 20 1820 80
rect 2680 20 2800 80
rect 1700 0 2800 20
rect 1700 -580 1720 0
rect 1780 -580 1800 0
rect 1700 -600 1800 -580
rect 2700 -20 2800 0
rect 2700 -600 2720 -20
rect 2780 -600 2800 -20
rect 1700 -620 2800 -600
rect 1700 -680 1820 -620
rect 2680 -680 2800 -620
rect 1700 -700 2800 -680
rect 5400 80 6500 100
rect 5400 20 5520 80
rect 6380 20 6500 80
rect 5400 0 6500 20
rect 5400 -20 5500 0
rect 5400 -580 5420 -20
rect 5480 -580 5500 -20
rect 5400 -600 5500 -580
rect 6400 -20 6500 0
rect 6400 -580 6420 -20
rect 6480 -580 6500 -20
rect 6400 -600 6500 -580
rect 5400 -620 6500 -600
rect 5400 -680 5520 -620
rect 6380 -680 6500 -620
rect 5400 -700 6500 -680
rect 2260 -847 6000 -840
rect 2260 -927 2380 -847
rect 5880 -927 6000 -847
rect 2260 -940 6000 -927
rect 2260 -965 2360 -940
rect 2260 -2242 2272 -965
rect 2348 -2242 2360 -965
rect 2260 -2250 2360 -2242
rect 5900 -962 6000 -940
rect 5900 -2239 5911 -962
rect 5987 -2239 6000 -962
rect 5900 -2250 6000 -2239
rect 2260 -2260 6000 -2250
rect 2260 -2340 2380 -2260
rect 5880 -2340 6000 -2260
rect 2260 -2350 6000 -2340
rect 1500 -2410 1600 -2380
rect 6600 -2380 6620 1880
rect 6680 -2380 6700 1880
rect 6600 -2410 6700 -2380
rect 1500 -2420 6700 -2410
rect 1500 -2500 1620 -2420
rect 6580 -2500 6700 -2420
rect 1500 -2510 6700 -2500
<< nsubdiff >>
rect -1600 3980 9800 4000
rect -1600 3820 -1380 3980
rect 9580 3820 9800 3980
rect -1600 3800 9800 3820
rect -1600 3780 -1400 3800
rect -1600 -4380 -1580 3780
rect -1420 -4380 -1400 3780
rect 9600 3780 9800 3800
rect -400 3680 8600 3700
rect -400 3620 -280 3680
rect 8480 3620 8600 3680
rect -400 3600 8600 3620
rect -400 3580 -300 3600
rect -400 2220 -380 3580
rect -320 2220 -300 3580
rect -400 2200 -300 2220
rect 8500 3580 8600 3600
rect 8500 2220 8520 3580
rect 8580 2220 8600 3580
rect 8500 2200 8600 2220
rect -400 2180 8600 2200
rect -400 2120 -280 2180
rect 8480 2120 8600 2180
rect -400 2100 8600 2120
rect -1000 1780 1000 1800
rect -1000 1720 -880 1780
rect 880 1720 1000 1780
rect -1000 1700 1000 1720
rect -1000 1680 -900 1700
rect -1000 320 -980 1680
rect -920 320 -900 1680
rect -1000 300 -900 320
rect 900 1680 1000 1700
rect 900 320 920 1680
rect 980 320 1000 1680
rect 900 300 1000 320
rect -1000 280 1000 300
rect -1000 220 -880 280
rect 880 220 1000 280
rect -1000 200 1000 220
rect -260 40 880 60
rect -260 -20 -140 40
rect 760 -20 880 40
rect -260 -40 880 -20
rect -260 -60 -160 -40
rect -260 -700 -240 -60
rect -180 -700 -160 -60
rect -260 -720 -160 -700
rect 780 -60 880 -40
rect 780 -700 800 -60
rect 860 -700 880 -60
rect 780 -720 880 -700
rect -260 -740 880 -720
rect -260 -800 -140 -740
rect 760 -800 880 -740
rect -260 -820 880 -800
rect -1300 -1020 1400 -1000
rect -1300 -1080 -1180 -1020
rect 1280 -1080 1400 -1020
rect -1300 -1100 1400 -1080
rect -1300 -1120 -1200 -1100
rect -1300 -2880 -1280 -1120
rect -1220 -2880 -1200 -1120
rect -1300 -2900 -1200 -2880
rect 1300 -1120 1400 -1100
rect 1300 -2880 1320 -1120
rect 1380 -2880 1400 -1120
rect 7200 1780 9200 1800
rect 7200 1720 7320 1780
rect 9080 1720 9200 1780
rect 7200 1700 9200 1720
rect 7200 1680 7300 1700
rect 7200 320 7220 1680
rect 7280 320 7300 1680
rect 7200 300 7300 320
rect 9100 1680 9200 1700
rect 9100 320 9120 1680
rect 9180 320 9200 1680
rect 9100 300 9200 320
rect 7200 280 9200 300
rect 7200 220 7320 280
rect 9080 220 9200 280
rect 7200 200 9200 220
rect 7320 60 8460 80
rect 7320 0 7440 60
rect 8340 0 8460 60
rect 7320 -20 8460 0
rect 7320 -40 7420 -20
rect 7320 -680 7340 -40
rect 7400 -680 7420 -40
rect 7320 -700 7420 -680
rect 8360 -40 8460 -20
rect 8360 -680 8380 -40
rect 8440 -680 8460 -40
rect 8360 -700 8460 -680
rect 7320 -720 8460 -700
rect 7320 -780 7440 -720
rect 8340 -780 8460 -720
rect 7320 -800 8460 -780
rect 6800 -1020 9500 -1000
rect 6800 -1080 6920 -1020
rect 9380 -1080 9500 -1020
rect 6800 -1100 9500 -1080
rect 6800 -1120 6900 -1100
rect 1300 -2900 1400 -2880
rect -1300 -2920 1400 -2900
rect -1300 -2980 -1180 -2920
rect 1280 -2980 1400 -2920
rect -1300 -3000 1400 -2980
rect 6800 -2880 6820 -1120
rect 6880 -2880 6900 -1120
rect 6800 -2900 6900 -2880
rect 9400 -1120 9500 -1100
rect 9400 -2880 9420 -1120
rect 9480 -2880 9500 -1120
rect 9400 -2900 9500 -2880
rect 6800 -2920 9500 -2900
rect 6800 -2980 6920 -2920
rect 9380 -2980 9500 -2920
rect 6800 -3000 9500 -2980
rect -700 -3120 900 -3100
rect -700 -3180 -580 -3120
rect 780 -3180 900 -3120
rect -700 -3200 900 -3180
rect -700 -3220 -600 -3200
rect -700 -4180 -680 -3220
rect -620 -4180 -600 -3220
rect -700 -4200 -600 -4180
rect 800 -3220 900 -3200
rect 800 -4180 820 -3220
rect 880 -4180 900 -3220
rect 800 -4200 900 -4180
rect -700 -4220 900 -4200
rect -700 -4280 -580 -4220
rect 780 -4280 900 -4220
rect -700 -4300 900 -4280
rect 7300 -3120 8900 -3100
rect 7300 -3180 7420 -3120
rect 8780 -3180 8900 -3120
rect 7300 -3200 8900 -3180
rect 7300 -3220 7400 -3200
rect 7300 -4180 7320 -3220
rect 7380 -4180 7400 -3220
rect 7300 -4200 7400 -4180
rect 8800 -3220 8900 -3200
rect 8800 -4180 8820 -3220
rect 8880 -4180 8900 -3220
rect 8800 -4200 8900 -4180
rect 7300 -4220 8900 -4200
rect 7300 -4280 7420 -4220
rect 8780 -4280 8900 -4220
rect 7300 -4300 8900 -4280
rect -1600 -4400 -1400 -4380
rect 9600 -4380 9620 3780
rect 9780 -4380 9800 3780
rect 9600 -4400 9800 -4380
rect -1600 -4420 9800 -4400
rect -1600 -4580 -1380 -4420
rect 9580 -4580 9800 -4420
rect -1600 -4600 9800 -4580
<< psubdiffcont >>
rect 1620 1920 6580 1980
rect 1520 -2380 1580 1880
rect 1820 1720 6380 1780
rect 1720 320 1780 1680
rect 6420 320 6480 1680
rect 1820 220 3040 280
rect 5160 220 6380 280
rect 1820 20 2680 80
rect 1720 -580 1780 0
rect 2720 -600 2780 -20
rect 1820 -680 2680 -620
rect 5520 20 6380 80
rect 5420 -580 5480 -20
rect 6420 -580 6480 -20
rect 5520 -680 6380 -620
rect 2380 -927 5880 -847
rect 2272 -2242 2348 -965
rect 5911 -2239 5987 -962
rect 2380 -2340 5880 -2260
rect 6620 -2380 6680 1880
rect 1620 -2500 6580 -2420
<< nsubdiffcont >>
rect -1380 3820 9580 3980
rect -1580 -4380 -1420 3780
rect -280 3620 8480 3680
rect -380 2220 -320 3580
rect 8520 2220 8580 3580
rect -280 2120 8480 2180
rect -880 1720 880 1780
rect -980 320 -920 1680
rect 920 320 980 1680
rect -880 220 880 280
rect -140 -20 760 40
rect -240 -700 -180 -60
rect 800 -700 860 -60
rect -140 -800 760 -740
rect -1180 -1080 1280 -1020
rect -1280 -2880 -1220 -1120
rect 1320 -2880 1380 -1120
rect 7320 1720 9080 1780
rect 7220 320 7280 1680
rect 9120 320 9180 1680
rect 7320 220 9080 280
rect 7440 0 8340 60
rect 7340 -680 7400 -40
rect 8380 -680 8440 -40
rect 7440 -780 8340 -720
rect 6920 -1080 9380 -1020
rect -1180 -2980 1280 -2920
rect 6820 -2880 6880 -1120
rect 9420 -2880 9480 -1120
rect 6920 -2980 9380 -2920
rect -580 -3180 780 -3120
rect -680 -4180 -620 -3220
rect 820 -4180 880 -3220
rect -580 -4280 780 -4220
rect 7420 -3180 8780 -3120
rect 7320 -4180 7380 -3220
rect 8820 -4180 8880 -3220
rect 7420 -4280 8780 -4220
rect 9620 -4380 9780 3780
rect -1380 -4580 9580 -4420
<< locali >>
rect -1600 3980 9800 4000
rect -1600 3920 -1580 3980
rect -1520 3920 -1480 3980
rect -1420 3920 -1380 3980
rect -1600 3880 -1380 3920
rect -1600 3820 -1580 3880
rect -1520 3820 -1480 3880
rect -1420 3820 -1380 3880
rect 9580 3820 9800 3980
rect -1600 3780 9800 3820
rect -1600 -4380 -1580 3780
rect -1420 3680 9620 3780
rect -1420 3620 -280 3680
rect 8480 3620 9620 3680
rect -1420 3600 9620 3620
rect -1420 3580 -300 3600
rect -1420 2220 -380 3580
rect -320 2220 -300 3580
rect 860 2400 980 3600
rect 2980 2400 3100 3600
rect 5100 2400 5220 3600
rect 7220 2400 7340 3600
rect 8500 3580 9620 3600
rect -1420 2200 -300 2220
rect 8500 2220 8520 3580
rect 8580 2220 9620 3580
rect 8500 2200 9620 2220
rect -1420 2180 9620 2200
rect -1420 2120 -280 2180
rect 8480 2120 9620 2180
rect -1420 2040 9620 2120
rect -1420 1780 1460 2040
rect -1420 1720 -880 1780
rect 880 1720 1460 1780
rect -1420 1700 1460 1720
rect -1420 1680 -900 1700
rect -1420 320 -980 1680
rect -920 320 -900 1680
rect 900 1680 1460 1700
rect -1420 300 -900 320
rect -440 300 -320 1440
rect 280 300 400 1440
rect 900 320 920 1680
rect 980 320 1460 1680
rect 900 300 1460 320
rect -1420 280 1460 300
rect -1420 220 -880 280
rect 880 220 1460 280
rect -1420 40 1460 220
rect -1420 -20 -140 40
rect 760 -20 1460 40
rect -1420 -40 1460 -20
rect -1420 -60 -160 -40
rect -1420 -700 -240 -60
rect -180 -340 -160 -60
rect 780 -60 1460 -40
rect -180 -420 260 -340
rect -180 -700 -160 -420
rect -1420 -720 -160 -700
rect 780 -700 800 -60
rect 860 -700 1460 -60
rect 780 -720 1460 -700
rect -1420 -740 1460 -720
rect -1420 -800 -140 -740
rect 760 -800 1460 -740
rect -1420 -1020 1460 -800
rect -1420 -1080 -1180 -1020
rect 1280 -1080 1460 -1020
rect -1420 -1100 1460 -1080
rect -1420 -1120 -1200 -1100
rect -1420 -2880 -1280 -1120
rect -1220 -2880 -1200 -1120
rect 1300 -1120 1460 -1100
rect -1420 -2900 -1200 -2880
rect -40 -2900 80 -1300
rect 1300 -2880 1320 -1120
rect 1380 -2560 1460 -1120
rect 1500 1980 6700 2000
rect 1500 1920 1620 1980
rect 6580 1920 6700 1980
rect 1500 1880 6700 1920
rect 1500 -2380 1520 1880
rect 1580 1780 6620 1880
rect 1580 1720 1820 1780
rect 6380 1720 6620 1780
rect 1580 1700 6620 1720
rect 1580 1680 1800 1700
rect 1580 320 1720 1680
rect 1780 320 1800 1680
rect 6400 1680 6620 1700
rect 1580 300 1800 320
rect 2940 300 3140 1440
rect 3720 440 3920 1340
rect 3720 380 3740 440
rect 3800 380 3840 440
rect 3900 380 3920 440
rect 3720 340 3920 380
rect 1580 280 3060 300
rect 1580 220 1820 280
rect 3040 220 3060 280
rect 3720 280 3740 340
rect 3800 280 3840 340
rect 3900 280 3920 340
rect 3720 260 3920 280
rect 4280 440 4480 1340
rect 4280 380 4300 440
rect 4360 380 4400 440
rect 4460 380 4480 440
rect 4280 340 4480 380
rect 4280 280 4300 340
rect 4360 280 4400 340
rect 4460 280 4480 340
rect 6400 320 6420 1680
rect 6480 320 6620 1680
rect 6400 300 6620 320
rect 4280 260 4480 280
rect 5140 280 6620 300
rect 1580 200 3060 220
rect 1580 80 3000 200
rect 3100 120 5100 260
rect 5140 220 5160 280
rect 6380 220 6620 280
rect 5140 200 6620 220
rect 1580 20 1820 80
rect 2680 20 3000 80
rect 1580 0 3000 20
rect 1580 -580 1720 0
rect 1780 -280 1800 0
rect 2700 -20 3000 0
rect 1780 -360 2240 -280
rect 1780 -580 1800 -360
rect 1580 -600 1800 -580
rect 2700 -600 2720 -20
rect 2780 -600 3000 -20
rect 1580 -620 3000 -600
rect 1580 -680 1820 -620
rect 2680 -680 3000 -620
rect 1580 -760 3000 -680
rect 5200 80 6620 200
rect 5200 20 5520 80
rect 6380 20 6620 80
rect 5200 0 6620 20
rect 5200 -20 5500 0
rect 5200 -580 5420 -20
rect 5480 -280 5500 -20
rect 6400 -20 6620 0
rect 5480 -360 5840 -280
rect 5480 -580 5500 -360
rect 5200 -600 5500 -580
rect 6400 -580 6420 -20
rect 6480 -580 6620 -20
rect 6400 -600 6620 -580
rect 5200 -620 6620 -600
rect 5200 -680 5520 -620
rect 6380 -680 6620 -620
rect 5200 -760 6620 -680
rect 1580 -847 6620 -760
rect 1580 -927 2380 -847
rect 5880 -927 6620 -847
rect 1580 -940 6620 -927
rect 1580 -965 2360 -940
rect 1580 -1080 2272 -965
rect 1580 -1140 1720 -1080
rect 1780 -1140 1980 -1080
rect 2040 -1140 2272 -1080
rect 1580 -1360 2272 -1140
rect 1580 -1420 1720 -1360
rect 1780 -1420 1980 -1360
rect 2040 -1420 2272 -1360
rect 1580 -2242 2272 -1420
rect 2348 -2242 2360 -965
rect 1580 -2250 2360 -2242
rect 5900 -962 6620 -940
rect 5900 -2239 5911 -962
rect 5987 -2239 6620 -962
rect 5900 -2250 6620 -2239
rect 1580 -2260 6620 -2250
rect 1580 -2340 2380 -2260
rect 5880 -2340 6620 -2260
rect 1580 -2380 6620 -2340
rect 6680 -2380 6700 1880
rect 1500 -2420 6700 -2380
rect 1500 -2500 1620 -2420
rect 6580 -2500 6700 -2420
rect 1500 -2510 6700 -2500
rect 6740 1780 9620 2040
rect 6740 1720 7320 1780
rect 9080 1720 9620 1780
rect 6740 1700 9620 1720
rect 6740 1680 7300 1700
rect 6740 320 7220 1680
rect 7280 320 7300 1680
rect 9100 1680 9620 1700
rect 6740 300 7300 320
rect 7760 300 7880 1440
rect 8480 300 8600 1440
rect 9100 320 9120 1680
rect 9180 320 9620 1680
rect 9100 300 9620 320
rect 6740 280 9620 300
rect 6740 220 7320 280
rect 9080 220 9620 280
rect 6740 60 9620 220
rect 6740 0 7440 60
rect 8340 0 9620 60
rect 6740 -20 9620 0
rect 6740 -40 7420 -20
rect 6740 -680 7340 -40
rect 7400 -680 7420 -40
rect 6740 -700 7420 -680
rect 7840 -700 7940 -20
rect 8360 -40 9620 -20
rect 8360 -680 8380 -40
rect 8440 -680 9620 -40
rect 8360 -700 9620 -680
rect 6740 -720 9620 -700
rect 6740 -780 7440 -720
rect 8340 -780 9620 -720
rect 6740 -1020 9620 -780
rect 6740 -1080 6920 -1020
rect 9380 -1080 9620 -1020
rect 6740 -1100 9620 -1080
rect 6740 -1120 6900 -1100
rect 6740 -2560 6820 -1120
rect 1380 -2880 6820 -2560
rect 6880 -2880 6900 -1120
rect 9400 -1120 9620 -1100
rect 1300 -2900 6900 -2880
rect 8060 -2900 8180 -1300
rect 9400 -2880 9420 -1120
rect 9480 -2880 9620 -1120
rect 9400 -2900 9620 -2880
rect -1420 -2920 9620 -2900
rect -1420 -2980 -1180 -2920
rect 1280 -2980 6920 -2920
rect 9380 -2980 9620 -2920
rect -1420 -3120 9620 -2980
rect -1420 -3180 -580 -3120
rect 780 -3180 7420 -3120
rect 8780 -3180 9620 -3120
rect -1420 -3200 9620 -3180
rect -1420 -3220 -600 -3200
rect -1420 -4180 -680 -3220
rect -620 -4180 -600 -3220
rect 800 -3220 7400 -3200
rect -1420 -4200 -600 -4180
rect -500 -4200 -380 -3400
rect 800 -4180 820 -3220
rect 880 -4180 7320 -3220
rect 7380 -4180 7400 -3220
rect 8800 -3220 9620 -3200
rect 800 -4200 7400 -4180
rect 8560 -4200 8680 -3400
rect 8800 -4180 8820 -3220
rect 8880 -4180 9620 -3220
rect 8800 -4200 9620 -4180
rect -1420 -4220 9620 -4200
rect -1420 -4280 -580 -4220
rect 780 -4280 7420 -4220
rect 8780 -4280 9620 -4220
rect -1420 -4380 9620 -4280
rect 9780 -4380 9800 3780
rect -1600 -4420 9800 -4380
rect -1600 -4580 -1380 -4420
rect 9580 -4580 9800 -4420
rect -1600 -4600 9800 -4580
<< viali >>
rect -1580 3920 -1520 3980
rect -1480 3920 -1420 3980
rect -1580 3820 -1520 3880
rect -1480 3820 -1420 3880
rect 3740 380 3800 440
rect 3840 380 3900 440
rect 3740 280 3800 340
rect 3840 280 3900 340
rect 4300 380 4360 440
rect 4400 380 4460 440
rect 4300 280 4360 340
rect 4400 280 4460 340
rect 1720 -1140 1780 -1080
rect 1980 -1140 2040 -1080
rect 1720 -1420 1780 -1360
rect 1980 -1420 2040 -1360
<< metal1 >>
rect -1600 3980 -1400 4000
rect -1600 3920 -1580 3980
rect -1520 3920 -1480 3980
rect -1420 3920 -1400 3980
rect -1600 3880 -1400 3920
rect -1600 3820 -1580 3880
rect -1520 3820 -1480 3880
rect -1420 3820 -1400 3880
rect -1600 3800 -1400 3820
rect -200 2980 0 3000
rect -200 2920 -180 2980
rect -120 2920 -80 2980
rect -20 2920 0 2980
rect -200 2880 0 2920
rect -200 2820 -180 2880
rect -120 2820 -80 2880
rect -20 2820 0 2880
rect -200 2800 0 2820
rect 1920 2360 2040 3400
rect 4000 2980 4200 3000
rect 4000 2920 4020 2980
rect 4080 2920 4120 2980
rect 4180 2920 4200 2980
rect 4000 2880 4200 2920
rect 4000 2820 4020 2880
rect 4080 2820 4120 2880
rect 4180 2820 4200 2880
rect 4000 2800 4200 2820
rect 6140 2360 6260 3400
rect 8220 2980 8420 3000
rect 8220 2920 8240 2980
rect 8300 2920 8340 2980
rect 8400 2920 8420 2980
rect 8220 2880 8420 2920
rect 8220 2820 8240 2880
rect 8300 2820 8340 2880
rect 8400 2820 8420 2880
rect 8220 2800 8420 2820
rect -100 2340 8240 2360
rect -100 2280 -80 2340
rect -20 2280 40 2340
rect 100 2280 160 2340
rect 220 2320 8240 2340
rect 220 2280 4060 2320
rect -100 2240 4060 2280
rect 4140 2240 8300 2320
rect -100 2200 8300 2240
rect -100 2180 4060 2200
rect -100 2120 -80 2180
rect -20 2120 40 2180
rect 100 2120 160 2180
rect 220 2120 4060 2180
rect 4140 2120 8300 2200
rect -100 2100 8300 2120
rect 820 1800 1100 2100
rect -700 1600 1100 1800
rect 7100 1800 7380 2100
rect 2380 1660 2580 1720
rect 2380 1620 2400 1660
rect -720 1500 1100 1600
rect 1940 1600 2400 1620
rect 2460 1600 2500 1660
rect 2560 1620 2580 1660
rect 5600 1660 5800 1720
rect 5600 1620 5620 1660
rect 2560 1600 5620 1620
rect 5680 1600 5720 1660
rect 5780 1620 5800 1660
rect 5780 1600 6240 1620
rect 1940 1560 6240 1600
rect 1940 1520 2400 1560
rect -800 300 -680 1440
rect -80 260 40 1440
rect 640 300 760 1440
rect 1940 1080 2060 1520
rect 2380 1500 2400 1520
rect 2460 1500 2500 1560
rect 2560 1520 5620 1560
rect 2560 1500 2580 1520
rect 2380 1480 2580 1500
rect 5600 1500 5620 1520
rect 5680 1500 5720 1560
rect 5780 1520 6240 1560
rect 5780 1500 5800 1520
rect 5600 1480 5800 1500
rect 1460 920 2060 1080
rect -800 140 760 260
rect -80 -160 40 140
rect -80 -200 340 -160
rect -80 -560 40 -200
rect 240 -240 340 -200
rect 1460 -300 1600 920
rect 1940 420 2060 920
rect 3720 1320 3920 1340
rect 3720 1260 3740 1320
rect 3800 1260 3840 1320
rect 3900 1260 3920 1320
rect 4280 1320 4480 1340
rect 3720 1220 3920 1260
rect 3720 1160 3740 1220
rect 3800 1160 3840 1220
rect 3900 1160 3920 1220
rect 3720 660 3920 1160
rect 3720 600 3740 660
rect 3800 600 3840 660
rect 3900 600 3920 660
rect 3720 560 3920 600
rect 3720 500 3740 560
rect 3800 500 3840 560
rect 3900 500 3920 560
rect 3720 440 3920 500
rect 4000 1220 4200 1300
rect 4000 1140 4060 1220
rect 4140 1140 4200 1220
rect 4000 1120 4200 1140
rect 4000 1040 4060 1120
rect 4140 1040 4200 1120
rect 4000 1020 4200 1040
rect 4000 940 4060 1020
rect 4140 940 4200 1020
rect 4000 920 4200 940
rect 4000 840 4060 920
rect 4140 840 4200 920
rect 4000 820 4200 840
rect 4000 740 4060 820
rect 4140 740 4200 820
rect 4000 720 4200 740
rect 4000 640 4060 720
rect 4140 640 4200 720
rect 4000 620 4200 640
rect 4000 540 4060 620
rect 4140 540 4200 620
rect 4000 520 4200 540
rect 4000 440 4060 520
rect 4140 440 4200 520
rect 4280 1260 4300 1320
rect 4360 1260 4400 1320
rect 4460 1260 4480 1320
rect 4280 1220 4480 1260
rect 4280 1160 4300 1220
rect 4360 1160 4400 1220
rect 4460 1160 4480 1220
rect 4280 660 4480 1160
rect 4280 600 4300 660
rect 4360 600 4400 660
rect 4460 600 4480 660
rect 4280 560 4480 600
rect 4280 500 4300 560
rect 4360 500 4400 560
rect 4460 500 4480 560
rect 4280 440 4480 500
rect 5060 1320 5260 1440
rect 5060 1260 5080 1320
rect 5140 1260 5180 1320
rect 5240 1260 5260 1320
rect 5060 1220 5260 1260
rect 5060 1160 5080 1220
rect 5140 1160 5180 1220
rect 5240 1160 5260 1220
rect 5060 660 5260 1160
rect 5060 600 5080 660
rect 5140 600 5180 660
rect 5240 600 5260 660
rect 5060 560 5260 600
rect 5060 500 5080 560
rect 5140 500 5180 560
rect 5240 500 5260 560
rect 5060 440 5260 500
rect 3720 380 3740 440
rect 3800 380 3840 440
rect 3900 380 3920 440
rect 3720 340 3920 380
rect 3720 280 3740 340
rect 3800 280 3840 340
rect 3900 280 3920 340
rect 3720 260 3920 280
rect 4280 380 4300 440
rect 4360 380 4400 440
rect 4460 380 4480 440
rect 6120 420 6240 1520
rect 7100 1500 8900 1800
rect 7400 1120 7520 1140
rect 7400 1040 7420 1120
rect 7500 1040 7520 1120
rect 7400 940 7520 1040
rect 7400 860 7420 940
rect 7500 860 7520 940
rect 7400 840 7520 860
rect 8120 1120 8240 1140
rect 8120 1040 8140 1120
rect 8220 1040 8240 1120
rect 8120 940 8240 1040
rect 8120 860 8140 940
rect 8220 860 8240 940
rect 8120 840 8240 860
rect 8840 1120 8960 1140
rect 8840 1040 8860 1120
rect 8940 1040 8960 1120
rect 8840 940 8960 1040
rect 8840 860 8860 940
rect 8940 860 8960 940
rect 8840 840 8960 860
rect 4280 340 4480 380
rect 4280 280 4300 340
rect 4360 280 4400 340
rect 4460 280 4480 340
rect 4280 260 4480 280
rect 6200 140 6400 160
rect 6200 80 6220 140
rect 6280 80 6320 140
rect 6380 80 6400 140
rect 6200 40 6400 80
rect 6200 -20 6220 40
rect 6280 -20 6320 40
rect 6380 -20 6400 40
rect 6200 -40 6400 -20
rect 340 -460 1600 -300
rect 1680 -120 2320 -100
rect 1680 -220 1700 -120
rect 1800 -220 1960 -120
rect 2060 -180 2320 -120
rect 5620 -180 5920 -100
rect 2060 -220 2080 -180
rect 1680 -400 2080 -220
rect 2300 -360 2720 -280
rect 1680 -500 1700 -400
rect 1800 -500 1960 -400
rect 2060 -440 2080 -400
rect 2060 -500 2320 -440
rect 1680 -520 2320 -500
rect 240 -560 340 -520
rect -80 -620 340 -560
rect 2640 -620 2720 -360
rect 5620 -440 5700 -180
rect 6260 -280 6340 -40
rect 7500 -120 8180 -40
rect 7500 -160 7580 -120
rect 5900 -360 6340 -280
rect 7220 -180 7580 -160
rect 7220 -260 7240 -180
rect 7320 -260 7380 -180
rect 7460 -260 7580 -180
rect 7220 -320 7580 -260
rect 7220 -400 7240 -320
rect 7320 -400 7380 -320
rect 7460 -400 7580 -320
rect 5620 -520 5920 -440
rect -80 -760 1540 -620
rect -1000 -940 1100 -900
rect -1000 -1020 840 -940
rect 920 -1020 980 -940
rect 1060 -1020 1100 -940
rect -1000 -1080 1100 -1020
rect -1000 -1140 840 -1080
rect -1020 -1160 840 -1140
rect 920 -1160 980 -1080
rect 1060 -1160 1100 -1080
rect -1020 -1240 1100 -1160
rect 1260 -1040 1540 -760
rect 2580 -640 2780 -620
rect 2580 -700 2600 -640
rect 2660 -700 2700 -640
rect 2760 -700 2780 -640
rect 2580 -740 2780 -700
rect 2580 -800 2600 -740
rect 2660 -800 2700 -740
rect 2760 -800 2780 -740
rect 2580 -820 2780 -800
rect 5820 -1040 5920 -520
rect 7220 -460 7580 -400
rect 7220 -540 7240 -460
rect 7320 -540 7380 -460
rect 7460 -540 7580 -460
rect 7220 -560 7580 -540
rect 8220 -560 9560 -160
rect 7500 -600 7580 -560
rect 7500 -680 8180 -600
rect 7100 -940 9200 -900
rect 7100 -1020 7160 -940
rect 7240 -1020 7300 -940
rect 7380 -1020 9200 -940
rect 1260 -1060 2740 -1040
rect 1260 -1160 1700 -1060
rect 1800 -1160 1960 -1060
rect 2060 -1160 2740 -1060
rect 1260 -1340 2740 -1160
rect 1260 -1440 1700 -1340
rect 1800 -1440 1960 -1340
rect 2060 -1440 2740 -1340
rect 1260 -1460 2740 -1440
rect 2800 -1480 3420 -1060
rect 3480 -1460 4100 -1040
rect 4160 -1460 4780 -1040
rect 4840 -1460 5460 -1040
rect 5520 -1060 6580 -1040
rect 5520 -1160 6040 -1060
rect 6140 -1160 6180 -1060
rect 6280 -1160 6320 -1060
rect 6420 -1160 6460 -1060
rect 6560 -1160 6580 -1060
rect 5520 -1200 6580 -1160
rect 7100 -1080 9200 -1020
rect 7100 -1160 7160 -1080
rect 7240 -1160 7300 -1080
rect 7380 -1160 9200 -1080
rect 7100 -1200 9200 -1160
rect 9260 -1060 9560 -560
rect 9260 -1160 9280 -1060
rect 9380 -1160 9440 -1060
rect 9540 -1160 9560 -1060
rect 9260 -1200 9560 -1160
rect 5520 -1300 6040 -1200
rect 6140 -1300 6180 -1200
rect 6280 -1300 6320 -1200
rect 6420 -1300 6460 -1200
rect 6560 -1300 6580 -1200
rect 7040 -1240 9160 -1200
rect 5520 -1340 6580 -1300
rect 5520 -1440 6040 -1340
rect 6140 -1440 6180 -1340
rect 6280 -1440 6320 -1340
rect 6420 -1440 6460 -1340
rect 6560 -1440 6580 -1340
rect 9260 -1300 9280 -1200
rect 9380 -1300 9440 -1200
rect 9540 -1300 9560 -1200
rect 9260 -1340 9560 -1300
rect 9260 -1440 9280 -1340
rect 9380 -1440 9440 -1340
rect 9540 -1440 9560 -1340
rect 5520 -1460 6580 -1440
rect -1080 -1880 -940 -1860
rect -1080 -1940 -1040 -1880
rect -980 -1940 -940 -1880
rect -1080 -1980 -940 -1940
rect -1080 -2040 -1040 -1980
rect -980 -2040 -940 -1980
rect -1080 -2080 -940 -2040
rect -1080 -2140 -1040 -2080
rect -980 -2140 -940 -2080
rect -1080 -2160 -940 -2140
rect 980 -1880 1120 -1860
rect 980 -1940 1020 -1880
rect 1080 -1940 1120 -1880
rect 980 -1980 1120 -1940
rect 980 -2040 1020 -1980
rect 1080 -2040 1120 -1980
rect 980 -2080 1120 -2040
rect 980 -2140 1020 -2080
rect 1080 -2140 1120 -2080
rect 980 -2160 1120 -2140
rect 2460 -2160 3080 -1740
rect 3140 -2140 3760 -1720
rect 3820 -2160 4440 -1740
rect 4500 -2160 5120 -1740
rect 5180 -2140 5800 -1720
rect 7000 -1880 7140 -1860
rect 7000 -1940 7040 -1880
rect 7100 -1940 7140 -1880
rect 7000 -1980 7140 -1940
rect 7000 -2040 7040 -1980
rect 7100 -2040 7140 -1980
rect 7000 -2080 7140 -2040
rect 7000 -2140 7040 -2080
rect 7100 -2140 7140 -2080
rect 7000 -2160 7140 -2140
rect 9060 -1880 9200 -1860
rect 9060 -1940 9100 -1880
rect 9160 -1940 9200 -1880
rect 9060 -1980 9200 -1940
rect 9060 -2040 9100 -1980
rect 9160 -2040 9200 -1980
rect 9060 -2080 9200 -2040
rect 9060 -2140 9100 -2080
rect 9160 -2140 9200 -2080
rect 9060 -2160 9200 -2140
rect -400 -3040 9260 -3020
rect -400 -3100 -380 -3040
rect -320 -3100 -260 -3040
rect -200 -3100 -140 -3040
rect -80 -3100 9260 -3040
rect -400 -3160 9260 -3100
rect -400 -3220 -380 -3160
rect -320 -3220 -260 -3160
rect -200 -3220 -140 -3160
rect -80 -3220 9260 -3160
rect -400 -3280 9260 -3220
rect -400 -3340 -380 -3280
rect -320 -3340 -260 -3280
rect -200 -3340 -140 -3280
rect -80 -3340 9260 -3280
rect -400 -3360 9260 -3340
rect 600 -3740 7600 -3720
rect 600 -3800 1140 -3740
rect 1200 -3800 1300 -3740
rect 1360 -3800 6840 -3740
rect 6900 -3800 7000 -3740
rect 7060 -3800 7600 -3740
rect 600 -3960 7600 -3800
rect 600 -4020 1140 -3960
rect 1200 -4020 1300 -3960
rect 1360 -4020 6840 -3960
rect 6900 -4020 7000 -3960
rect 7060 -4020 7600 -3960
rect 600 -4040 7600 -4020
<< via1 >>
rect -180 2920 -120 2980
rect -80 2920 -20 2980
rect -180 2820 -120 2880
rect -80 2820 -20 2880
rect 4020 2920 4080 2980
rect 4120 2920 4180 2980
rect 4020 2820 4080 2880
rect 4120 2820 4180 2880
rect 8240 2920 8300 2980
rect 8340 2920 8400 2980
rect 8240 2820 8300 2880
rect 8340 2820 8400 2880
rect -80 2280 -20 2340
rect 40 2280 100 2340
rect 160 2280 220 2340
rect 4060 2240 4140 2320
rect -80 2120 -20 2180
rect 40 2120 100 2180
rect 160 2120 220 2180
rect 4060 2120 4140 2200
rect 2400 1600 2460 1660
rect 2500 1600 2560 1660
rect 5620 1600 5680 1660
rect 5720 1600 5780 1660
rect 2400 1500 2460 1560
rect 2500 1500 2560 1560
rect 5620 1500 5680 1560
rect 5720 1500 5780 1560
rect 3740 1260 3800 1320
rect 3840 1260 3900 1320
rect 3740 1160 3800 1220
rect 3840 1160 3900 1220
rect 3740 600 3800 660
rect 3840 600 3900 660
rect 3740 500 3800 560
rect 3840 500 3900 560
rect 4060 1140 4140 1220
rect 4060 1040 4140 1120
rect 4060 940 4140 1020
rect 4060 840 4140 920
rect 4060 740 4140 820
rect 4060 640 4140 720
rect 4060 540 4140 620
rect 4060 440 4140 520
rect 4300 1260 4360 1320
rect 4400 1260 4460 1320
rect 4300 1160 4360 1220
rect 4400 1160 4460 1220
rect 4300 600 4360 660
rect 4400 600 4460 660
rect 4300 500 4360 560
rect 4400 500 4460 560
rect 5080 1260 5140 1320
rect 5180 1260 5240 1320
rect 5080 1160 5140 1220
rect 5180 1160 5240 1220
rect 5080 600 5140 660
rect 5180 600 5240 660
rect 5080 500 5140 560
rect 5180 500 5240 560
rect 7420 1040 7500 1120
rect 7420 860 7500 940
rect 8140 1040 8220 1120
rect 8140 860 8220 940
rect 8860 1040 8940 1120
rect 8860 860 8940 940
rect 6220 80 6280 140
rect 6320 80 6380 140
rect 6220 -20 6280 40
rect 6320 -20 6380 40
rect 1700 -220 1800 -120
rect 1960 -220 2060 -120
rect 1700 -500 1800 -400
rect 1960 -500 2060 -400
rect 7240 -260 7320 -180
rect 7380 -260 7460 -180
rect 7240 -400 7320 -320
rect 7380 -400 7460 -320
rect 840 -1020 920 -940
rect 980 -1020 1060 -940
rect 840 -1160 920 -1080
rect 980 -1160 1060 -1080
rect 2600 -700 2660 -640
rect 2700 -700 2760 -640
rect 2600 -800 2660 -740
rect 2700 -800 2760 -740
rect 7240 -540 7320 -460
rect 7380 -540 7460 -460
rect 7160 -1020 7240 -940
rect 7300 -1020 7380 -940
rect 1700 -1080 1800 -1060
rect 1700 -1140 1720 -1080
rect 1720 -1140 1780 -1080
rect 1780 -1140 1800 -1080
rect 1700 -1160 1800 -1140
rect 1960 -1080 2060 -1060
rect 1960 -1140 1980 -1080
rect 1980 -1140 2040 -1080
rect 2040 -1140 2060 -1080
rect 1960 -1160 2060 -1140
rect 1700 -1360 1800 -1340
rect 1700 -1420 1720 -1360
rect 1720 -1420 1780 -1360
rect 1780 -1420 1800 -1360
rect 1700 -1440 1800 -1420
rect 1960 -1360 2060 -1340
rect 1960 -1420 1980 -1360
rect 1980 -1420 2040 -1360
rect 2040 -1420 2060 -1360
rect 1960 -1440 2060 -1420
rect 6040 -1160 6140 -1060
rect 6180 -1160 6280 -1060
rect 6320 -1160 6420 -1060
rect 6460 -1160 6560 -1060
rect 7160 -1160 7240 -1080
rect 7300 -1160 7380 -1080
rect 9280 -1160 9380 -1060
rect 9440 -1160 9540 -1060
rect 6040 -1300 6140 -1200
rect 6180 -1300 6280 -1200
rect 6320 -1300 6420 -1200
rect 6460 -1300 6560 -1200
rect 6040 -1440 6140 -1340
rect 6180 -1440 6280 -1340
rect 6320 -1440 6420 -1340
rect 6460 -1440 6560 -1340
rect 9280 -1300 9380 -1200
rect 9440 -1300 9540 -1200
rect 9280 -1440 9380 -1340
rect 9440 -1440 9540 -1340
rect -1040 -1940 -980 -1880
rect -1040 -2040 -980 -1980
rect -1040 -2140 -980 -2080
rect 1020 -1940 1080 -1880
rect 1020 -2040 1080 -1980
rect 1020 -2140 1080 -2080
rect 7040 -1940 7100 -1880
rect 7040 -2040 7100 -1980
rect 7040 -2140 7100 -2080
rect 9100 -1940 9160 -1880
rect 9100 -2040 9160 -1980
rect 9100 -2140 9160 -2080
rect -380 -3100 -320 -3040
rect -260 -3100 -200 -3040
rect -140 -3100 -80 -3040
rect -380 -3220 -320 -3160
rect -260 -3220 -200 -3160
rect -140 -3220 -80 -3160
rect -380 -3340 -320 -3280
rect -260 -3340 -200 -3280
rect -140 -3340 -80 -3280
rect 1140 -3800 1200 -3740
rect 1300 -3800 1360 -3740
rect 6840 -3800 6900 -3740
rect 7000 -3800 7060 -3740
rect 1140 -4020 1200 -3960
rect 1300 -4020 1360 -3960
rect 6840 -4020 6900 -3960
rect 7000 -4020 7060 -3960
<< metal2 >>
rect -180 2980 8420 3000
rect -120 2920 -80 2980
rect -20 2920 4020 2980
rect 4080 2920 4120 2980
rect 4180 2920 8240 2980
rect 8300 2920 8340 2980
rect 8400 2920 8420 2980
rect -180 2880 8420 2920
rect -120 2820 -80 2880
rect -20 2820 4020 2880
rect 4080 2820 4120 2880
rect 4180 2820 8240 2880
rect 8300 2820 8340 2880
rect 8400 2820 8420 2880
rect -180 2800 8420 2820
rect -1480 2340 240 2360
rect -1480 2280 -1460 2340
rect -1400 2280 -1340 2340
rect -1280 2280 -1220 2340
rect -1160 2280 -80 2340
rect -20 2280 40 2340
rect 100 2280 160 2340
rect 220 2280 240 2340
rect -1480 2180 240 2280
rect -1480 2120 -1460 2180
rect -1400 2120 -1340 2180
rect -1280 2120 -1220 2180
rect -1160 2120 -80 2180
rect -20 2120 40 2180
rect 100 2120 160 2180
rect 220 2120 240 2180
rect -1480 2100 240 2120
rect 2380 1660 2580 2800
rect 2380 1600 2400 1660
rect 2460 1600 2500 1660
rect 2560 1600 2580 1660
rect 2380 1560 2580 1600
rect 2380 1500 2400 1560
rect 2460 1500 2500 1560
rect 2560 1500 2580 1560
rect 2380 1480 2580 1500
rect 4000 2320 4200 2360
rect 4000 2240 4060 2320
rect 4140 2240 4200 2320
rect 4000 2200 4200 2240
rect 4000 2120 4060 2200
rect 4140 2120 4200 2200
rect 3720 1320 3920 1340
rect 3720 1260 3740 1320
rect 3800 1260 3840 1320
rect 3900 1260 3920 1320
rect 3720 1220 3920 1260
rect 3720 1160 3740 1220
rect 3800 1160 3840 1220
rect 3900 1160 3920 1220
rect 3720 1140 3920 1160
rect 4000 1220 4200 2120
rect 5600 1660 5800 2800
rect 5600 1600 5620 1660
rect 5680 1600 5720 1660
rect 5780 1600 5800 1660
rect 5600 1560 5800 1600
rect 5600 1500 5620 1560
rect 5680 1500 5720 1560
rect 5780 1500 5800 1560
rect 5600 1480 5800 1500
rect 4000 1140 4060 1220
rect 4140 1140 4200 1220
rect 4280 1320 4480 1340
rect 4280 1260 4300 1320
rect 4360 1260 4400 1320
rect 4460 1260 4480 1320
rect 4280 1220 4480 1260
rect 4280 1160 4300 1220
rect 4360 1160 4400 1220
rect 4460 1160 4480 1220
rect 4280 1140 4480 1160
rect 5060 1320 5260 1340
rect 5060 1260 5080 1320
rect 5140 1260 5180 1320
rect 5240 1260 5260 1320
rect 5060 1220 5260 1260
rect 5060 1160 5080 1220
rect 5140 1160 5180 1220
rect 5240 1160 5260 1220
rect 5060 1140 5260 1160
rect 4000 1120 4200 1140
rect 4000 1040 4060 1120
rect 4140 1040 4200 1120
rect 4000 1020 4200 1040
rect 4000 940 4060 1020
rect 4140 940 4200 1020
rect 4000 920 4200 940
rect 4000 840 4060 920
rect 4140 840 4200 920
rect 4000 820 4200 840
rect 4000 740 4060 820
rect 4140 740 4200 820
rect 4000 720 4200 740
rect 3720 660 3920 680
rect 3720 600 3740 660
rect 3800 600 3840 660
rect 3900 600 3920 660
rect 3720 560 3920 600
rect 3720 500 3740 560
rect 3800 500 3840 560
rect 3900 500 3920 560
rect 3720 480 3920 500
rect 4000 640 4060 720
rect 4140 640 4200 720
rect 7200 1120 9200 1140
rect 7200 1040 7420 1120
rect 7500 1040 8140 1120
rect 8220 1040 8860 1120
rect 8940 1040 9200 1120
rect 7200 940 9200 1040
rect 7200 860 7420 940
rect 7500 860 8140 940
rect 8220 860 8860 940
rect 8940 860 9200 940
rect 7200 840 9200 860
rect 4000 620 4200 640
rect 4000 540 4060 620
rect 4140 540 4200 620
rect 4000 520 4200 540
rect 4000 440 4060 520
rect 4140 440 4200 520
rect 4280 660 4480 680
rect 4280 600 4300 660
rect 4360 600 4400 660
rect 4460 600 4480 660
rect 4280 560 4480 600
rect 4280 500 4300 560
rect 4360 500 4400 560
rect 4460 500 4480 560
rect 4280 480 4480 500
rect 5060 660 5260 680
rect 5060 600 5080 660
rect 5140 600 5180 660
rect 5240 600 5260 660
rect 5060 560 5260 600
rect 5060 500 5080 560
rect 5140 500 5180 560
rect 5240 500 5260 560
rect 5060 480 5260 500
rect 4000 400 4200 440
rect 7200 160 7480 840
rect 1680 140 7480 160
rect 1680 80 6220 140
rect 6280 80 6320 140
rect 6380 80 7480 140
rect 1680 40 7480 80
rect 1680 -20 6220 40
rect 6280 -20 6320 40
rect 6380 -20 7480 40
rect 1680 -40 7480 -20
rect 1680 -120 2080 -40
rect 1680 -220 1700 -120
rect 1800 -220 1960 -120
rect 2060 -220 2080 -120
rect 1680 -400 2080 -220
rect 1680 -500 1700 -400
rect 1800 -500 1960 -400
rect 2060 -500 2080 -400
rect 820 -940 1080 -920
rect 820 -1020 840 -940
rect 920 -1020 980 -940
rect 1060 -1020 1080 -940
rect 820 -1080 1080 -1020
rect 820 -1160 840 -1080
rect 920 -1160 980 -1080
rect 1060 -1160 1080 -1080
rect 820 -1180 1080 -1160
rect 1680 -1060 2080 -500
rect 7220 -180 7480 -160
rect 7220 -260 7240 -180
rect 7320 -260 7380 -180
rect 7460 -260 7480 -180
rect 7220 -320 7480 -260
rect 7220 -400 7240 -320
rect 7320 -400 7380 -320
rect 7460 -400 7480 -320
rect 7220 -460 7480 -400
rect 7220 -540 7240 -460
rect 7320 -540 7380 -460
rect 7460 -540 7480 -460
rect 7220 -620 7480 -540
rect 2440 -640 7480 -620
rect 2440 -700 2600 -640
rect 2660 -700 2700 -640
rect 2760 -700 7480 -640
rect 2440 -740 7480 -700
rect 2440 -800 2600 -740
rect 2660 -800 2700 -740
rect 2760 -800 7480 -740
rect 2440 -820 7480 -800
rect 7140 -940 7400 -820
rect 7140 -1020 7160 -940
rect 7240 -1020 7300 -940
rect 7380 -1020 7400 -940
rect 1680 -1160 1700 -1060
rect 1800 -1160 1960 -1060
rect 2060 -1160 2080 -1060
rect 1680 -1340 2080 -1160
rect 1680 -1440 1700 -1340
rect 1800 -1440 1960 -1340
rect 2060 -1440 2080 -1340
rect 1680 -1460 2080 -1440
rect 6020 -1060 6580 -1040
rect 6020 -1160 6040 -1060
rect 6140 -1160 6180 -1060
rect 6280 -1160 6320 -1060
rect 6420 -1160 6460 -1060
rect 6560 -1160 6580 -1060
rect 6020 -1200 6580 -1160
rect 7140 -1080 7400 -1020
rect 7140 -1160 7160 -1080
rect 7240 -1160 7300 -1080
rect 7380 -1160 7400 -1080
rect 7140 -1180 7400 -1160
rect 9260 -1060 9560 -1040
rect 9260 -1160 9280 -1060
rect 9380 -1160 9440 -1060
rect 9540 -1160 9560 -1060
rect 6020 -1300 6040 -1200
rect 6140 -1300 6180 -1200
rect 6280 -1300 6320 -1200
rect 6420 -1300 6460 -1200
rect 6560 -1220 6580 -1200
rect 9260 -1200 9560 -1160
rect 9260 -1220 9280 -1200
rect 6560 -1300 9280 -1220
rect 9380 -1300 9440 -1200
rect 9540 -1300 9560 -1200
rect 6020 -1340 9560 -1300
rect 6020 -1440 6040 -1340
rect 6140 -1440 6180 -1340
rect 6280 -1440 6320 -1340
rect 6420 -1440 6460 -1340
rect 6560 -1420 9280 -1340
rect 6560 -1440 6580 -1420
rect 6020 -1460 6580 -1440
rect 9260 -1440 9280 -1420
rect 9380 -1440 9440 -1340
rect 9540 -1440 9560 -1340
rect 9260 -1460 9560 -1440
rect -1080 -1880 1380 -1860
rect -1080 -1940 -1040 -1880
rect -980 -1940 1020 -1880
rect 1080 -1940 1380 -1880
rect -1080 -1980 1380 -1940
rect -1080 -2040 -1040 -1980
rect -980 -2040 1020 -1980
rect 1080 -2040 1380 -1980
rect -1080 -2080 1380 -2040
rect -1080 -2140 -1040 -2080
rect -980 -2140 1020 -2080
rect 1080 -2140 1380 -2080
rect -1080 -2160 1380 -2140
rect -1480 -3040 -60 -3020
rect -1480 -3100 -1460 -3040
rect -1400 -3100 -1340 -3040
rect -1280 -3100 -1220 -3040
rect -1160 -3100 -380 -3040
rect -320 -3100 -260 -3040
rect -200 -3100 -140 -3040
rect -80 -3100 -60 -3040
rect -1480 -3160 -60 -3100
rect -1480 -3220 -1460 -3160
rect -1400 -3220 -1340 -3160
rect -1280 -3220 -1220 -3160
rect -1160 -3220 -380 -3160
rect -320 -3220 -260 -3160
rect -200 -3220 -140 -3160
rect -80 -3220 -60 -3160
rect -1480 -3280 -60 -3220
rect -1480 -3340 -1460 -3280
rect -1400 -3340 -1340 -3280
rect -1280 -3340 -1220 -3280
rect -1160 -3340 -380 -3280
rect -320 -3340 -260 -3280
rect -200 -3340 -140 -3280
rect -80 -3340 -60 -3280
rect -1480 -3360 -60 -3340
rect 1120 -3740 1380 -2160
rect 1120 -3800 1140 -3740
rect 1200 -3800 1300 -3740
rect 1360 -3800 1380 -3740
rect 1120 -3960 1380 -3800
rect 1120 -4020 1140 -3960
rect 1200 -4020 1300 -3960
rect 1360 -4020 1380 -3960
rect 1120 -4040 1380 -4020
rect 6820 -1880 9200 -1860
rect 6820 -1940 7040 -1880
rect 7100 -1940 9100 -1880
rect 9160 -1940 9200 -1880
rect 6820 -1980 9200 -1940
rect 6820 -2040 7040 -1980
rect 7100 -2040 9100 -1980
rect 9160 -2040 9200 -1980
rect 6820 -2080 9200 -2040
rect 6820 -2140 7040 -2080
rect 7100 -2140 9100 -2080
rect 9160 -2140 9200 -2080
rect 6820 -2160 9200 -2140
rect 6820 -3740 7080 -2160
rect 6820 -3800 6840 -3740
rect 6900 -3800 7000 -3740
rect 7060 -3800 7080 -3740
rect 6820 -3960 7080 -3800
rect 6820 -4020 6840 -3960
rect 6900 -4020 7000 -3960
rect 7060 -4020 7080 -3960
rect 6820 -4040 7080 -4020
<< via2 >>
rect -1460 2280 -1400 2340
rect -1340 2280 -1280 2340
rect -1220 2280 -1160 2340
rect -1460 2120 -1400 2180
rect -1340 2120 -1280 2180
rect -1220 2120 -1160 2180
rect 3740 1260 3800 1320
rect 3840 1260 3900 1320
rect 3740 1160 3800 1220
rect 3840 1160 3900 1220
rect 4300 1260 4360 1320
rect 4400 1260 4460 1320
rect 4300 1160 4360 1220
rect 4400 1160 4460 1220
rect 5080 1260 5140 1320
rect 5180 1260 5240 1320
rect 5080 1160 5140 1220
rect 5180 1160 5240 1220
rect 3740 600 3800 660
rect 3840 600 3900 660
rect 3740 500 3800 560
rect 3840 500 3900 560
rect 4300 600 4360 660
rect 4400 600 4460 660
rect 4300 500 4360 560
rect 4400 500 4460 560
rect 5080 600 5140 660
rect 5180 600 5240 660
rect 5080 500 5140 560
rect 5180 500 5240 560
rect 840 -1000 900 -940
rect 1000 -1000 1060 -940
rect 840 -1160 900 -1100
rect 1000 -1160 1060 -1100
rect 7160 -1000 7220 -940
rect 7320 -1000 7380 -940
rect 7160 -1160 7220 -1100
rect 7320 -1160 7380 -1100
rect -1460 -3100 -1400 -3040
rect -1340 -3100 -1280 -3040
rect -1220 -3100 -1160 -3040
rect -1460 -3220 -1400 -3160
rect -1340 -3220 -1280 -3160
rect -1220 -3220 -1160 -3160
rect -1460 -3340 -1400 -3280
rect -1340 -3340 -1280 -3280
rect -1220 -3340 -1160 -3280
<< metal3 >>
rect -1480 2340 -1140 2360
rect -1480 2280 -1460 2340
rect -1400 2280 -1340 2340
rect -1280 2280 -1220 2340
rect -1160 2280 -1140 2340
rect -1480 2180 -1140 2280
rect -1480 2120 -1460 2180
rect -1400 2120 -1340 2180
rect -1280 2120 -1220 2180
rect -1160 2120 -1140 2180
rect -1480 -3040 -1140 2120
rect 3720 1320 5260 1340
rect 3720 1260 3740 1320
rect 3800 1260 3840 1320
rect 3900 1260 4300 1320
rect 4360 1260 4400 1320
rect 4460 1260 5080 1320
rect 5140 1260 5180 1320
rect 5240 1260 5260 1320
rect 3720 1220 5260 1260
rect 3720 1160 3740 1220
rect 3800 1160 3840 1220
rect 3900 1160 4300 1220
rect 4360 1160 4400 1220
rect 4460 1160 5080 1220
rect 5140 1160 5180 1220
rect 5240 1160 5260 1220
rect 3720 1140 5260 1160
rect 3720 660 5260 680
rect 3720 600 3740 660
rect 3800 600 3840 660
rect 3900 600 4300 660
rect 4360 600 4400 660
rect 4460 600 5080 660
rect 5140 600 5180 660
rect 5240 600 5260 660
rect 3720 560 5260 600
rect 3720 500 3740 560
rect 3800 500 3840 560
rect 3900 500 4300 560
rect 4360 500 4400 560
rect 4460 500 5080 560
rect 5140 500 5180 560
rect 5240 500 5260 560
rect 3720 480 5260 500
rect 800 -940 7440 -900
rect 800 -1000 840 -940
rect 900 -1000 1000 -940
rect 1060 -1000 7160 -940
rect 7220 -1000 7320 -940
rect 7380 -1000 7440 -940
rect 800 -1100 7440 -1000
rect 800 -1160 840 -1100
rect 900 -1160 1000 -1100
rect 1060 -1160 7160 -1100
rect 7220 -1160 7320 -1100
rect 7380 -1160 7440 -1100
rect 800 -1240 7440 -1160
rect -1480 -3100 -1460 -3040
rect -1400 -3100 -1340 -3040
rect -1280 -3100 -1220 -3040
rect -1160 -3100 -1140 -3040
rect -1480 -3160 -1140 -3100
rect -1480 -3220 -1460 -3160
rect -1400 -3220 -1340 -3160
rect -1280 -3220 -1220 -3160
rect -1160 -3220 -1140 -3160
rect -1480 -3280 -1140 -3220
rect -1480 -3340 -1460 -3280
rect -1400 -3340 -1340 -3280
rect -1280 -3340 -1220 -3280
rect -1160 -3340 -1140 -3280
rect -1480 -3360 -1140 -3340
use sky130_fd_pr__res_generic_l1_58A49Y  R1
timestamp 1770979109
transform 1 0 3400 0 1 -333
box -100 -467 100 467
use sky130_fd_pr__res_generic_l1_58A49Y  R3
timestamp 1770979109
transform 1 0 3600 0 1 -333
box -100 -467 100 467
use sky130_fd_pr__res_generic_l1_58A49Y  R4
timestamp 1770979109
transform 1 0 3800 0 1 -333
box -100 -467 100 467
use sky130_fd_pr__res_generic_l1_58A49Y  R5
timestamp 1770979109
transform 1 0 4000 0 1 -333
box -100 -467 100 467
use sky130_fd_pr__res_generic_l1_58A49Y  R6
timestamp 1770979109
transform 1 0 4200 0 1 -333
box -100 -467 100 467
use sky130_fd_pr__res_generic_l1_58A49Y  R7
timestamp 1770979109
transform 1 0 4400 0 1 -333
box -100 -467 100 467
use sky130_fd_pr__res_generic_l1_58A49Y  R8
timestamp 1770979109
transform 1 0 4600 0 1 -333
box -100 -467 100 467
use sky130_fd_pr__res_generic_l1_58A49Y  R9
timestamp 1770979109
transform 1 0 4800 0 1 -333
box -100 -467 100 467
use sky130_fd_pr__res_generic_l1_58A49Y  R10
timestamp 1770979109
transform 1 0 5000 0 1 -333
box -100 -467 100 467
use sky130_fd_pr__res_generic_l1_58A49Y  R21
timestamp 1770979109
transform 1 0 3200 0 1 -333
box -100 -467 100 467
use sky130_fd_pr__nfet_01v8_RX9YJP  sky130_fd_pr__nfet_01v8_RX9YJP_0
timestamp 1770979109
transform 1 0 5873 0 1 -312
box -73 -188 73 188
use sky130_fd_pr__pfet_01v8_AW5DE3  sky130_fd_pr__pfet_01v8_AW5DE3_0
timestamp 1770979109
transform 1 0 8181 0 1 998
box -781 -598 781 564
use sky130_fd_pr__pfet_01v8_MW3DW6  sky130_fd_pr__pfet_01v8_MW3DW6_0
timestamp 1770979109
transform 1 0 8123 0 1 -1977
box -1123 -823 1123 789
use sky130_fd_pr__pfet_01v8_VCUNPM  sky130_fd_pr__pfet_01v8_VCUNPM_0
timestamp 1770979109
transform 1 0 8094 0 1 -3689
box -594 -411 594 377
use sky130_fd_pr__res_xhigh_po_1p41_CGMGNJ  sky130_fd_pr__res_xhigh_po_1p41_CGMGNJ_0
timestamp 1770979109
transform 1 0 2601 0 1 -1593
box -141 -557 141 557
use sky130_fd_pr__nfet_01v8_CEKAWC  XM1
timestamp 1770979109
transform 1 0 4098 0 1 1010
box -2145 -557 2145 557
use sky130_fd_pr__pfet_01v8_WYTN36  XM3
timestamp 1770979109
transform 1 0 4097 0 1 2864
box -4297 -564 4297 598
use sky130_fd_pr__pfet_01v8_Y44983  XM5
timestamp 1770979109
transform 1 0 289 0 1 -380
box -109 -200 109 200
use sky130_fd_pr__pfet_01v8_AW5DE3  XM6
timestamp 1770979109
transform 1 0 -19 0 1 998
box -781 -598 781 564
use sky130_fd_pr__pfet_01v8_FX5EQP  XM8
timestamp 1770979109
transform 1 0 7883 0 1 -360
box -423 -300 423 300
use sky130_fd_pr__pfet_01v8_VCUNPM  XM10
timestamp 1770979109
transform 1 0 94 0 1 -3689
box -594 -411 594 377
use sky130_fd_pr__pfet_01v8_MW3DW6  XM11
timestamp 1770979109
transform 1 0 23 0 1 -1977
box -1123 -823 1123 789
use sky130_fd_pr__nfet_01v8_RX9YJP  XM13
timestamp 1770979109
transform 1 0 2273 0 1 -312
box -73 -188 73 188
use sky130_fd_pr__res_xhigh_po_1p41_CGMGNJ  XR2
timestamp 1770979109
transform 1 0 2941 0 1 -1593
box -141 -557 141 557
use sky130_fd_pr__res_xhigh_po_1p41_CGMGNJ  XR12
timestamp 1770979109
transform 1 0 3281 0 1 -1593
box -141 -557 141 557
use sky130_fd_pr__res_xhigh_po_1p41_CGMGNJ  XR13
timestamp 1770979109
transform 1 0 3621 0 1 -1593
box -141 -557 141 557
use sky130_fd_pr__res_xhigh_po_1p41_CGMGNJ  XR14
timestamp 1770979109
transform 1 0 3961 0 1 -1593
box -141 -557 141 557
use sky130_fd_pr__res_xhigh_po_1p41_CGMGNJ  XR15
timestamp 1770979109
transform 1 0 4301 0 1 -1593
box -141 -557 141 557
use sky130_fd_pr__res_xhigh_po_1p41_CGMGNJ  XR16
timestamp 1770979109
transform 1 0 4641 0 1 -1593
box -141 -557 141 557
use sky130_fd_pr__res_xhigh_po_1p41_CGMGNJ  XR17
timestamp 1770979109
transform 1 0 4981 0 1 -1593
box -141 -557 141 557
use sky130_fd_pr__res_xhigh_po_1p41_CGMGNJ  XR18
timestamp 1770979109
transform 1 0 5321 0 1 -1593
box -141 -557 141 557
use sky130_fd_pr__res_xhigh_po_1p41_CGMGNJ  XR19
timestamp 1770979109
transform 1 0 5661 0 1 -1593
box -141 -557 141 557
<< labels >>
flabel metal1 -1600 3800 -1400 4000 0 FreeSans 1600 0 0 0 VDD
port 4 nsew
flabel metal1 1360 -4040 6840 -3720 0 FreeSans 1600 0 0 0 IREF
port 6 nsew
flabel locali 1580 -2420 2272 -1420 0 FreeSans 1600 0 0 0 VSS
port 8 nsew
<< end >>

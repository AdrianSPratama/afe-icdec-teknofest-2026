magic
tech sky130A
magscale 1 10
timestamp 1771420802
<< error_p >>
rect 24760 44430 33940 44490
rect 24760 14800 24820 44430
rect 24940 44250 33760 44310
rect 24940 43730 25000 44250
rect 25005 43730 25085 43810
rect 25155 43730 25235 43810
rect 33465 43730 33545 43810
rect 33615 43730 33695 43810
rect 33700 43730 33760 44250
rect 24925 43650 25005 43730
rect 25235 43650 25315 43730
rect 33385 43650 33465 43730
rect 33695 43650 33775 43730
rect 24940 14800 25000 43650
rect 25695 42212 25775 42292
rect 25845 42212 25925 42292
rect 27465 42212 27545 42292
rect 27615 42212 27695 42292
rect 29235 42212 29315 42292
rect 29385 42212 29465 42292
rect 31005 42212 31085 42292
rect 31155 42212 31235 42292
rect 32775 42212 32855 42292
rect 32925 42212 33005 42292
rect 25615 42132 25695 42212
rect 25925 42132 26005 42212
rect 27385 42132 27465 42212
rect 27695 42132 27775 42212
rect 29155 42132 29235 42212
rect 29465 42132 29545 42212
rect 30925 42132 31005 42212
rect 31235 42132 31315 42212
rect 32695 42132 32775 42212
rect 33005 42132 33085 42212
rect 25615 39528 25695 39608
rect 25925 39528 26005 39608
rect 27385 39528 27465 39608
rect 27695 39528 27775 39608
rect 29155 39528 29235 39608
rect 29465 39528 29545 39608
rect 30925 39528 31005 39608
rect 31235 39528 31315 39608
rect 32695 39528 32775 39608
rect 33005 39528 33085 39608
rect 25695 39448 25775 39528
rect 25845 39448 25925 39528
rect 27465 39448 27545 39528
rect 27615 39448 27695 39528
rect 29235 39448 29315 39528
rect 29385 39448 29465 39528
rect 31005 39448 31085 39528
rect 31155 39448 31235 39528
rect 32775 39448 32855 39528
rect 32925 39448 33005 39528
rect 26345 38120 27045 38190
rect 28115 38120 28815 38190
rect 29885 38120 30585 38190
rect 31655 38120 32355 38190
rect 26580 37955 26660 38035
rect 26730 37955 26810 38035
rect 28350 37955 28430 38035
rect 28500 37955 28580 38035
rect 30120 37955 30200 38035
rect 30270 37955 30350 38035
rect 31890 37955 31970 38035
rect 32040 37955 32120 38035
rect 26500 37875 26890 37955
rect 28270 37875 28660 37955
rect 30040 37875 30430 37955
rect 31810 37875 32200 37955
rect 26525 37805 26865 37875
rect 28295 37805 28635 37875
rect 30065 37805 30405 37875
rect 31835 37805 32175 37875
rect 26500 37725 26890 37805
rect 28270 37725 28660 37805
rect 30040 37725 30430 37805
rect 31810 37725 32200 37805
rect 26580 37645 26660 37725
rect 26730 37645 26810 37725
rect 28350 37645 28430 37725
rect 28500 37645 28580 37725
rect 30120 37645 30200 37725
rect 30270 37645 30350 37725
rect 31890 37645 31970 37725
rect 32040 37645 32120 37725
rect 25695 35792 25775 35872
rect 25845 35792 25925 35872
rect 27465 35792 27545 35872
rect 27615 35792 27695 35872
rect 29235 35792 29315 35872
rect 29385 35792 29465 35872
rect 31005 35792 31085 35872
rect 31155 35792 31235 35872
rect 32775 35792 32855 35872
rect 32925 35792 33005 35872
rect 25615 35712 25695 35792
rect 25925 35712 26005 35792
rect 27385 35712 27465 35792
rect 27695 35712 27775 35792
rect 29155 35712 29235 35792
rect 29465 35712 29545 35792
rect 30925 35712 31005 35792
rect 31235 35712 31315 35792
rect 32695 35712 32775 35792
rect 33005 35712 33085 35792
rect 25615 33108 25695 33188
rect 25925 33108 26005 33188
rect 27385 33108 27465 33188
rect 27695 33108 27775 33188
rect 29155 33108 29235 33188
rect 29465 33108 29545 33188
rect 30925 33108 31005 33188
rect 31235 33108 31315 33188
rect 32695 33108 32775 33188
rect 33005 33108 33085 33188
rect 25695 33028 25775 33108
rect 25845 33028 25925 33108
rect 27465 33028 27545 33108
rect 27615 33028 27695 33108
rect 29235 33028 29315 33108
rect 29385 33028 29465 33108
rect 31005 33028 31085 33108
rect 31155 33028 31235 33108
rect 32775 33028 32855 33108
rect 32925 33028 33005 33108
rect 26345 31700 27045 31770
rect 28115 31700 28815 31770
rect 29885 31700 30585 31770
rect 31655 31700 32355 31770
rect 26580 31535 26660 31615
rect 26730 31535 26810 31615
rect 28350 31535 28430 31615
rect 28500 31535 28580 31615
rect 30120 31535 30200 31615
rect 30270 31535 30350 31615
rect 31890 31535 31970 31615
rect 32040 31535 32120 31615
rect 26500 31455 26890 31535
rect 28270 31455 28660 31535
rect 30040 31455 30430 31535
rect 31810 31455 32200 31535
rect 26525 31385 26865 31455
rect 28295 31385 28635 31455
rect 30065 31385 30405 31455
rect 31835 31385 32175 31455
rect 26500 31305 26890 31385
rect 28270 31305 28660 31385
rect 30040 31305 30430 31385
rect 31810 31305 32200 31385
rect 26580 31225 26660 31305
rect 26730 31225 26810 31305
rect 28350 31225 28430 31305
rect 28500 31225 28580 31305
rect 30120 31225 30200 31305
rect 30270 31225 30350 31305
rect 31890 31225 31970 31305
rect 32040 31225 32120 31305
rect 25695 29372 25775 29452
rect 25845 29372 25925 29452
rect 27465 29372 27545 29452
rect 27615 29372 27695 29452
rect 29235 29372 29315 29452
rect 29385 29372 29465 29452
rect 31005 29372 31085 29452
rect 31155 29372 31235 29452
rect 32775 29372 32855 29452
rect 32925 29372 33005 29452
rect 25615 29292 25695 29372
rect 25925 29292 26005 29372
rect 27385 29292 27465 29372
rect 27695 29292 27775 29372
rect 29155 29292 29235 29372
rect 29465 29292 29545 29372
rect 30925 29292 31005 29372
rect 31235 29292 31315 29372
rect 32695 29292 32775 29372
rect 33005 29292 33085 29372
rect 25615 26688 25695 26768
rect 25925 26688 26005 26768
rect 27385 26688 27465 26768
rect 27695 26688 27775 26768
rect 29155 26688 29235 26768
rect 29465 26688 29545 26768
rect 30925 26688 31005 26768
rect 31235 26688 31315 26768
rect 32695 26688 32775 26768
rect 33005 26688 33085 26768
rect 25695 26608 25775 26688
rect 25845 26608 25925 26688
rect 27465 26608 27545 26688
rect 27615 26608 27695 26688
rect 29235 26608 29315 26688
rect 29385 26608 29465 26688
rect 31005 26608 31085 26688
rect 31155 26608 31235 26688
rect 32775 26608 32855 26688
rect 32925 26608 33005 26688
rect 26345 25280 27045 25350
rect 28115 25280 28815 25350
rect 29885 25280 30585 25350
rect 31655 25280 32355 25350
rect 26580 25115 26660 25195
rect 26730 25115 26810 25195
rect 28350 25115 28430 25195
rect 28500 25115 28580 25195
rect 30120 25115 30200 25195
rect 30270 25115 30350 25195
rect 31890 25115 31970 25195
rect 32040 25115 32120 25195
rect 26500 25035 26890 25115
rect 28270 25035 28660 25115
rect 30040 25035 30430 25115
rect 31810 25035 32200 25115
rect 26525 24965 26865 25035
rect 28295 24965 28635 25035
rect 30065 24965 30405 25035
rect 31835 24965 32175 25035
rect 26500 24885 26890 24965
rect 28270 24885 28660 24965
rect 30040 24885 30430 24965
rect 31810 24885 32200 24965
rect 26580 24805 26660 24885
rect 26730 24805 26810 24885
rect 28350 24805 28430 24885
rect 28500 24805 28580 24885
rect 30120 24805 30200 24885
rect 30270 24805 30350 24885
rect 31890 24805 31970 24885
rect 32040 24805 32120 24885
rect 25695 22952 25775 23032
rect 25845 22952 25925 23032
rect 27465 22952 27545 23032
rect 27615 22952 27695 23032
rect 29235 22952 29315 23032
rect 29385 22952 29465 23032
rect 31005 22952 31085 23032
rect 31155 22952 31235 23032
rect 32775 22952 32855 23032
rect 32925 22952 33005 23032
rect 25615 22872 25695 22952
rect 25925 22872 26005 22952
rect 27385 22872 27465 22952
rect 27695 22872 27775 22952
rect 29155 22872 29235 22952
rect 29465 22872 29545 22952
rect 30925 22872 31005 22952
rect 31235 22872 31315 22952
rect 32695 22872 32775 22952
rect 33005 22872 33085 22952
rect 25615 20268 25695 20348
rect 25925 20268 26005 20348
rect 27385 20268 27465 20348
rect 27695 20268 27775 20348
rect 29155 20268 29235 20348
rect 29465 20268 29545 20348
rect 30925 20268 31005 20348
rect 31235 20268 31315 20348
rect 32695 20268 32775 20348
rect 33005 20268 33085 20348
rect 25695 20188 25775 20268
rect 25845 20188 25925 20268
rect 27465 20188 27545 20268
rect 27615 20188 27695 20268
rect 29235 20188 29315 20268
rect 29385 20188 29465 20268
rect 31005 20188 31085 20268
rect 31155 20188 31235 20268
rect 32775 20188 32855 20268
rect 32925 20188 33005 20268
rect 26345 18860 27045 18930
rect 28115 18860 28815 18930
rect 29885 18860 30585 18930
rect 31655 18860 32355 18930
rect 26580 18695 26660 18775
rect 26730 18695 26810 18775
rect 28350 18695 28430 18775
rect 28500 18695 28580 18775
rect 30120 18695 30200 18775
rect 30270 18695 30350 18775
rect 31890 18695 31970 18775
rect 32040 18695 32120 18775
rect 26500 18615 26890 18695
rect 28270 18615 28660 18695
rect 30040 18615 30430 18695
rect 31810 18615 32200 18695
rect 26525 18545 26865 18615
rect 28295 18545 28635 18615
rect 30065 18545 30405 18615
rect 31835 18545 32175 18615
rect 26500 18465 26890 18545
rect 28270 18465 28660 18545
rect 30040 18465 30430 18545
rect 31810 18465 32200 18545
rect 26580 18385 26660 18465
rect 26730 18385 26810 18465
rect 28350 18385 28430 18465
rect 28500 18385 28580 18465
rect 30120 18385 30200 18465
rect 30270 18385 30350 18465
rect 31890 18385 31970 18465
rect 32040 18385 32120 18465
rect 25695 16532 25775 16612
rect 25845 16532 25925 16612
rect 27465 16532 27545 16612
rect 27615 16532 27695 16612
rect 29235 16532 29315 16612
rect 29385 16532 29465 16612
rect 31005 16532 31085 16612
rect 31155 16532 31235 16612
rect 32775 16532 32855 16612
rect 32925 16532 33005 16612
rect 25615 16452 25695 16532
rect 25925 16452 26005 16532
rect 27385 16452 27465 16532
rect 27695 16452 27775 16532
rect 29155 16452 29235 16532
rect 29465 16452 29545 16532
rect 30925 16452 31005 16532
rect 31235 16452 31315 16532
rect 32695 16452 32775 16532
rect 33005 16452 33085 16532
rect 33700 14800 33760 43650
rect 33880 14800 33940 44430
<< error_s >>
rect 24760 11390 24820 14800
rect 24940 12170 25000 14800
rect 25615 13848 25695 13928
rect 25925 13848 26005 13928
rect 27385 13848 27465 13928
rect 27695 13848 27775 13928
rect 29155 13848 29235 13928
rect 29465 13848 29545 13928
rect 30925 13848 31005 13928
rect 31235 13848 31315 13928
rect 32695 13848 32775 13928
rect 33005 13848 33085 13928
rect 25695 13768 25775 13848
rect 25845 13768 25925 13848
rect 27465 13768 27545 13848
rect 27615 13768 27695 13848
rect 29235 13768 29315 13848
rect 29385 13768 29465 13848
rect 31005 13768 31085 13848
rect 31155 13768 31235 13848
rect 32775 13768 32855 13848
rect 32925 13768 33005 13848
rect 26345 12440 27045 12510
rect 28115 12440 28815 12510
rect 29885 12440 30585 12510
rect 31655 12440 32355 12510
rect 26580 12275 26660 12355
rect 26730 12275 26810 12355
rect 28350 12275 28430 12355
rect 28500 12275 28580 12355
rect 30120 12275 30200 12355
rect 30270 12275 30350 12355
rect 31890 12275 31970 12355
rect 32040 12275 32120 12355
rect 26500 12195 26890 12275
rect 28270 12195 28660 12275
rect 30040 12195 30430 12275
rect 31810 12195 32200 12275
rect 24925 12090 25005 12170
rect 25235 12090 25315 12170
rect 26525 12125 26865 12195
rect 28295 12125 28635 12195
rect 30065 12125 30405 12195
rect 31835 12125 32175 12195
rect 33700 12170 33760 14800
rect 24940 11570 25000 12090
rect 25005 12010 25085 12090
rect 25155 12010 25235 12090
rect 26500 12045 26890 12125
rect 28270 12045 28660 12125
rect 30040 12045 30430 12125
rect 31810 12045 32200 12125
rect 33385 12090 33465 12170
rect 33695 12090 33775 12170
rect 26580 11965 26660 12045
rect 26730 11965 26810 12045
rect 28350 11965 28430 12045
rect 28500 11965 28580 12045
rect 30120 11965 30200 12045
rect 30270 11965 30350 12045
rect 31890 11965 31970 12045
rect 32040 11965 32120 12045
rect 33465 12010 33545 12090
rect 33615 12010 33695 12090
rect 33700 11570 33760 12090
rect 24940 11510 33760 11570
rect 33880 11390 33940 14800
rect 24760 11330 33940 11390
rect 6795 -1450 7085 -1420
rect 17295 -1450 17585 -1420
rect 6795 -1620 6855 -1450
rect 17295 -1620 17355 -1450
rect 6795 -1650 7085 -1620
rect 17295 -1650 17585 -1620
rect -10420 -3590 -10400 -3080
rect 13390 -3200 13400 -3050
rect 13530 -3060 13540 -2910
rect -10280 -3450 -10260 -3220
rect 10295 -3250 10585 -3220
rect 13795 -3250 14085 -3220
rect 10295 -3420 10355 -3250
rect 13795 -3420 13855 -3250
rect 10295 -3450 10585 -3420
rect 13795 -3450 14085 -3420
rect -4900 -4600 -4790 -4580
rect -5040 -4770 -4960 -4750
rect 10295 -5950 10585 -5920
rect 13795 -5950 14085 -5920
rect 10295 -6120 10355 -5950
rect 13795 -6120 13855 -5950
rect 10295 -6150 10585 -6120
rect 13795 -6150 14085 -6120
rect 6700 -6200 6900 -6170
rect 7000 -6200 7200 -6170
rect 6560 -6340 6760 -6310
rect 7120 -6340 7340 -6310
rect 13390 -6350 13400 -6170
rect 17200 -6200 17400 -6170
rect 17480 -6200 17700 -6170
rect 13530 -6490 13540 -6310
rect 17060 -6340 17260 -6310
rect 17620 -6340 17840 -6310
rect 6795 -7750 7085 -7720
rect 17295 -7750 17585 -7720
rect 6795 -7920 6855 -7750
rect 17295 -7920 17355 -7750
rect 6795 -7950 7085 -7920
rect 17295 -7950 17585 -7920
<< nwell >>
rect -12200 700 29700 7200
rect 20300 -27200 29700 700
<< pwell >>
rect -12000 -17000 20000 500
<< psubdiff >>
rect -7500 400 -500 500
rect -7500 100 -6900 400
rect -1100 100 -500 400
rect -7500 0 -500 100
rect -7500 -100 -7000 0
rect -12000 -600 -8000 -500
rect -12000 -900 -11400 -600
rect -8600 -900 -8000 -600
rect -12000 -1000 -8000 -900
rect -12000 -1100 -11500 -1000
rect -12000 -3900 -11900 -1100
rect -11600 -3900 -11500 -1100
rect -12000 -4000 -11500 -3900
rect -8500 -1100 -8000 -1000
rect -8500 -3900 -8400 -1100
rect -8100 -3900 -8000 -1100
rect -8500 -4000 -8000 -3900
rect -12000 -4100 -8000 -4000
rect -12000 -4400 -11400 -4100
rect -8600 -4400 -8000 -4100
rect -12000 -4500 -8000 -4400
rect -7500 -5400 -7400 -100
rect -7100 -5400 -7000 -100
rect -7500 -5500 -7000 -5400
rect -1000 -100 -500 0
rect -1000 -5400 -900 -100
rect -600 -5400 -500 -100
rect -1000 -5500 -500 -5400
rect -7500 -5600 -500 -5500
rect -7500 -5900 -6900 -5600
rect -1100 -5900 -500 -5600
rect -7500 -6000 -500 -5900
rect 4500 400 20000 500
rect 4500 100 5100 400
rect 19400 100 20000 400
rect 4500 0 20000 100
rect 4500 -100 5000 0
rect -12000 -6600 -2500 -6500
rect -12000 -6900 -11400 -6600
rect -3100 -6900 -2500 -6600
rect -12000 -7000 -2500 -6900
rect -12000 -7100 -11500 -7000
rect -12000 -16400 -11900 -7100
rect -11600 -16400 -11500 -7100
rect -12000 -16500 -11500 -16400
rect -3000 -7100 -2500 -7000
rect -3000 -16400 -2900 -7100
rect -2600 -16400 -2500 -7100
rect 4500 -9400 4600 -100
rect 4900 -9400 5000 -100
rect 19500 -100 20000 0
rect 5500 -600 8500 -500
rect 5500 -900 5800 -600
rect 8200 -900 8500 -600
rect 5500 -1000 8500 -900
rect 5500 -4000 6000 -1000
rect 8000 -4000 8500 -1000
rect 5500 -4500 8500 -4000
rect 9000 -600 12000 -500
rect 9000 -900 9300 -600
rect 11700 -900 12000 -600
rect 9000 -1000 12000 -900
rect 9000 -4000 9500 -1000
rect 11500 -4000 12000 -1000
rect 9000 -4500 12000 -4000
rect 12500 -600 15500 -500
rect 12500 -900 12800 -600
rect 15200 -900 15500 -600
rect 12500 -1000 15500 -900
rect 12500 -4000 13000 -1000
rect 15000 -4000 15500 -1000
rect 12500 -4500 15500 -4000
rect 16000 -600 19000 -500
rect 16000 -900 16300 -600
rect 18700 -900 19000 -600
rect 16000 -1000 19000 -900
rect 16000 -4000 16500 -1000
rect 18500 -4000 19000 -1000
rect 16000 -4500 19000 -4000
rect 5500 -5500 8500 -5000
rect 5500 -8500 6000 -5500
rect 8000 -8500 8500 -5500
rect 5500 -8600 8500 -8500
rect 5500 -8900 5800 -8600
rect 8200 -8900 8500 -8600
rect 5500 -9000 8500 -8900
rect 9000 -5500 12000 -5000
rect 9000 -8500 9500 -5500
rect 11500 -8500 12000 -5500
rect 9000 -8600 12000 -8500
rect 9000 -8900 9300 -8600
rect 11700 -8900 12000 -8600
rect 9000 -9000 12000 -8900
rect 12500 -5500 15500 -5000
rect 12500 -8500 13000 -5500
rect 15000 -8500 15500 -5500
rect 12500 -8600 15500 -8500
rect 12500 -8900 12800 -8600
rect 15200 -8900 15500 -8600
rect 12500 -9000 15500 -8900
rect 16000 -5500 19000 -5000
rect 16000 -8500 16500 -5500
rect 18500 -8500 19000 -5500
rect 16000 -8600 19000 -8500
rect 16000 -8900 16300 -8600
rect 18700 -8900 19000 -8600
rect 16000 -9000 19000 -8900
rect 4500 -9500 5000 -9400
rect 19500 -9400 19600 -100
rect 19900 -9400 20000 -100
rect 19500 -9500 20000 -9400
rect 4500 -9600 20000 -9500
rect 4500 -9900 5100 -9600
rect 19400 -9900 20000 -9600
rect 4500 -10000 20000 -9900
rect -3000 -16500 -2500 -16400
rect 4500 -10600 8500 -10500
rect 4500 -10900 5000 -10600
rect 8000 -10900 8500 -10600
rect 4500 -11000 8500 -10900
rect 4500 -11100 5000 -11000
rect 4500 -15900 4600 -11100
rect 4900 -15900 5000 -11100
rect 4500 -16000 5000 -15900
rect 8000 -11100 8500 -11000
rect 8000 -15900 8100 -11100
rect 8400 -15900 8500 -11100
rect 8000 -16000 8500 -15900
rect 4500 -16100 8500 -16000
rect 4500 -16400 5000 -16100
rect 8000 -16400 8500 -16100
rect 4500 -16500 8500 -16400
rect 11500 -10600 20000 -10500
rect 11500 -10900 12100 -10600
rect 19400 -10900 20000 -10600
rect 11500 -11000 20000 -10900
rect 11500 -11100 12000 -11000
rect 11500 -15900 11600 -11100
rect 11900 -15900 12000 -11100
rect 11500 -16000 12000 -15900
rect 19500 -11100 20000 -11000
rect 19500 -15900 19600 -11100
rect 19900 -15900 20000 -11100
rect 19500 -16000 20000 -15900
rect 11500 -16100 20000 -16000
rect 11500 -16400 12100 -16100
rect 19400 -16400 20000 -16100
rect 11500 -16500 20000 -16400
rect -12000 -16600 -2500 -16500
rect -12000 -16900 -11400 -16600
rect -3100 -16900 -2500 -16600
rect -12000 -17000 -2500 -16900
<< nsubdiff >>
rect -12000 6900 4000 7000
rect -12000 6600 -11400 6900
rect 3400 6600 4000 6900
rect -12000 6500 4000 6600
rect -12000 6400 -11500 6500
rect -12000 1600 -11900 6400
rect -11600 1600 -11500 6400
rect -12000 1500 -11500 1600
rect 3500 6400 4000 6500
rect 3500 1600 3600 6400
rect 3900 1600 4000 6400
rect 3500 1500 4000 1600
rect -12000 1400 4000 1500
rect -12000 1100 -11400 1400
rect 3400 1100 4000 1400
rect -12000 1000 4000 1100
rect 4500 6900 20000 7000
rect 4500 6600 5100 6900
rect 19400 6600 20000 6900
rect 4500 6500 20000 6600
rect 4500 6400 5000 6500
rect 4500 1600 4600 6400
rect 4900 1600 5000 6400
rect 4500 1500 5000 1600
rect 19500 6400 20000 6500
rect 19500 1600 19600 6400
rect 19900 1600 20000 6400
rect 19500 1500 20000 1600
rect 4500 1400 20000 1500
rect 4500 1100 5100 1400
rect 19400 1100 20000 1400
rect 4500 1000 20000 1100
rect 20500 6900 29500 7000
rect 20500 6600 21100 6900
rect 28900 6600 29500 6900
rect 20500 6500 29500 6600
rect 20500 6400 21000 6500
rect 20500 -26400 20600 6400
rect 20900 -26400 21000 6400
rect 20500 -26500 21000 -26400
rect 29000 6400 29500 6500
rect 29000 -26400 29100 6400
rect 29400 -26400 29500 6400
rect 29000 -26500 29500 -26400
rect 20500 -26600 29500 -26500
rect 20500 -26900 21100 -26600
rect 28900 -26900 29500 -26600
rect 20500 -27000 29500 -26900
<< psubdiffcont >>
rect -6900 100 -1100 400
rect -11400 -900 -8600 -600
rect -11900 -3900 -11600 -1100
rect -8400 -3900 -8100 -1100
rect -11400 -4400 -8600 -4100
rect -7400 -5400 -7100 -100
rect -900 -5400 -600 -100
rect -6900 -5900 -1100 -5600
rect 5100 100 19400 400
rect -11400 -6900 -3100 -6600
rect -11900 -16400 -11600 -7100
rect -2900 -16400 -2600 -7100
rect 4600 -9400 4900 -100
rect 5800 -900 8200 -600
rect 9300 -900 11700 -600
rect 12800 -900 15200 -600
rect 16300 -900 18700 -600
rect 5800 -8900 8200 -8600
rect 9300 -8900 11700 -8600
rect 12800 -8900 15200 -8600
rect 16300 -8900 18700 -8600
rect 19600 -9400 19900 -100
rect 5100 -9900 19400 -9600
rect 5000 -10900 8000 -10600
rect 4600 -15900 4900 -11100
rect 8100 -15900 8400 -11100
rect 5000 -16400 8000 -16100
rect 12100 -10900 19400 -10600
rect 11600 -15900 11900 -11100
rect 19600 -15900 19900 -11100
rect 12100 -16400 19400 -16100
rect -11400 -16900 -3100 -16600
<< nsubdiffcont >>
rect -11400 6600 3400 6900
rect -11900 1600 -11600 6400
rect 3600 1600 3900 6400
rect -11400 1100 3400 1400
rect 5100 6600 19400 6900
rect 4600 1600 4900 6400
rect 19600 1600 19900 6400
rect 5100 1100 19400 1400
rect 21100 6600 28900 6900
rect 20600 -26400 20900 6400
rect 29100 -26400 29400 6400
rect 21100 -26900 28900 -26600
<< locali >>
rect -12000 10400 -2500 10500
rect -12000 10100 -11900 10400
rect -11600 10100 -2500 10400
rect -12000 9900 -2500 10100
rect -12000 9600 -11900 9900
rect -11600 9600 -2500 9900
rect -12000 9400 -2500 9600
rect -12000 9100 -11900 9400
rect -11600 9100 -2500 9400
rect -12000 8900 -2500 9100
rect -12000 8600 -11900 8900
rect -11600 8600 -2500 8900
rect -12000 8400 -2500 8600
rect -12000 8100 -11900 8400
rect -11600 8100 -2500 8400
rect -12000 7900 -2500 8100
rect -12000 7600 -11900 7900
rect -11600 7600 -2500 7900
rect -12000 7400 -2500 7600
rect -12000 7100 -11900 7400
rect -11600 7100 -2500 7400
rect -12000 7000 -2500 7100
rect -12000 6900 4000 7000
rect -12000 6600 -11400 6900
rect 3400 6600 4000 6900
rect -12000 6500 4000 6600
rect -12000 6400 -11500 6500
rect -12000 1600 -11900 6400
rect -11600 1600 -11500 6400
rect -9400 2600 -8900 6500
rect -6300 2600 -5800 6500
rect -2400 2600 -1900 6500
rect 700 2600 1200 6500
rect 3500 6400 4000 6500
rect -12000 1500 -11500 1600
rect 3500 1600 3600 6400
rect 3900 1600 4000 6400
rect 3500 1500 4000 1600
rect -12000 1400 4000 1500
rect -12000 1100 -11400 1400
rect 3400 1100 4000 1400
rect -12000 1000 4000 1100
rect 4500 6900 20000 7000
rect 4500 6600 5100 6900
rect 19400 6600 20000 6900
rect 4500 6500 20000 6600
rect 4500 6400 5000 6500
rect 4500 1600 4600 6400
rect 4900 1600 5000 6400
rect 7500 3000 8000 6500
rect 10500 3000 11000 6500
rect 13500 3000 14000 6500
rect 16500 3000 17000 6500
rect 19500 6400 20000 6500
rect 4500 1500 5000 1600
rect 19500 1600 19600 6400
rect 19900 1600 20000 6400
rect 19500 1500 20000 1600
rect 4500 1400 20000 1500
rect 4500 1100 5100 1400
rect 19400 1100 20000 1400
rect 4500 1000 20000 1100
rect 20500 6900 29500 7000
rect 20500 6600 21100 6900
rect 28900 6600 29500 6900
rect 20500 6500 29500 6600
rect 20500 6400 21000 6500
rect -7500 400 -500 500
rect -7500 100 -6900 400
rect -1100 100 -500 400
rect -7500 0 -500 100
rect -7500 -100 -7000 0
rect -12000 -600 -8000 -500
rect -12000 -900 -11400 -600
rect -8600 -900 -8000 -600
rect -12000 -1000 -8000 -900
rect -12000 -1100 -11500 -1000
rect -12000 -3900 -11900 -1100
rect -11600 -3900 -11500 -1100
rect -12000 -4000 -11500 -3900
rect -8500 -1100 -8000 -1000
rect -8500 -3900 -8400 -1100
rect -8100 -3900 -8000 -1100
rect -8500 -4000 -8000 -3900
rect -12000 -4100 -8000 -4000
rect -12000 -4400 -11400 -4100
rect -8600 -4400 -8000 -4100
rect -12000 -4500 -8000 -4400
rect -7500 -5400 -7400 -100
rect -7100 -5400 -7000 -100
rect -4900 -4600 -4400 0
rect -1000 -100 -500 0
rect -7500 -5500 -7000 -5400
rect -1000 -5400 -900 -100
rect -600 -5400 -500 -100
rect -1000 -5500 -500 -5400
rect -7500 -5600 -500 -5500
rect -7500 -5900 -6900 -5600
rect -1100 -5900 -500 -5600
rect -7500 -6000 -500 -5900
rect 4500 400 20000 500
rect 4500 100 5100 400
rect 19400 100 20000 400
rect 4500 -100 20000 100
rect -12000 -6600 -2500 -6500
rect -12000 -6900 -11400 -6600
rect -3100 -6900 -2500 -6600
rect -12000 -7000 -2500 -6900
rect -12000 -7100 -11500 -7000
rect -12000 -16400 -11900 -7100
rect -11600 -16400 -11500 -7100
rect -12000 -16500 -11500 -16400
rect -3000 -7100 -2500 -7000
rect -3000 -16400 -2900 -7100
rect -2600 -16400 -2500 -7100
rect 4500 -9400 4600 -100
rect 4900 -300 19600 -100
rect 4900 -9200 5300 -300
rect 5700 -600 8300 -500
rect 5700 -900 5800 -600
rect 8200 -900 8300 -600
rect 5700 -1000 8300 -900
rect 8500 -4500 9000 -500
rect 9200 -600 11800 -500
rect 9200 -900 9300 -600
rect 11700 -900 11800 -600
rect 9200 -1000 11800 -900
rect 12000 -600 12500 -500
rect 12000 -900 12100 -600
rect 12400 -900 12500 -600
rect 12000 -1100 12500 -900
rect 12700 -600 15300 -500
rect 12700 -900 12800 -600
rect 15200 -900 15300 -600
rect 12700 -1000 15300 -900
rect 12000 -1400 12100 -1100
rect 12400 -1400 12500 -1100
rect 12000 -1600 12500 -1400
rect 12000 -1900 12100 -1600
rect 12400 -1900 12500 -1600
rect 12000 -2100 12500 -1900
rect 12000 -2400 12100 -2100
rect 12400 -2400 12500 -2100
rect 12000 -2600 12500 -2400
rect 12000 -2900 12100 -2600
rect 12400 -2900 12500 -2600
rect 12000 -3100 12500 -2900
rect 12000 -3400 12100 -3100
rect 12400 -3400 12500 -3100
rect 12000 -4500 12500 -3400
rect 15500 -4500 16000 -500
rect 16200 -600 18800 -500
rect 16200 -900 16300 -600
rect 18700 -900 18800 -600
rect 16200 -1000 18800 -900
rect 5500 -5000 19000 -4500
rect 5700 -8600 8300 -8500
rect 5700 -8900 5800 -8600
rect 8200 -8900 8300 -8600
rect 5700 -9000 8300 -8900
rect 8500 -9000 9000 -5000
rect 12000 -6100 12500 -5000
rect 12000 -6400 12100 -6100
rect 12400 -6400 12500 -6100
rect 12000 -6600 12500 -6400
rect 12000 -6900 12100 -6600
rect 12400 -6900 12500 -6600
rect 12000 -7100 12500 -6900
rect 12000 -7400 12100 -7100
rect 12400 -7400 12500 -7100
rect 12000 -7600 12500 -7400
rect 12000 -7900 12100 -7600
rect 12400 -7900 12500 -7600
rect 12000 -8100 12500 -7900
rect 12000 -8400 12100 -8100
rect 12400 -8400 12500 -8100
rect 9200 -8600 11800 -8500
rect 9200 -8900 9300 -8600
rect 11700 -8900 11800 -8600
rect 9200 -9000 11800 -8900
rect 12000 -8600 12500 -8400
rect 12000 -8900 12100 -8600
rect 12400 -8900 12500 -8600
rect 12000 -9000 12500 -8900
rect 12700 -8600 15300 -8500
rect 12700 -8900 12800 -8600
rect 15200 -8900 15300 -8600
rect 12700 -9000 15300 -8900
rect 15500 -9000 16000 -5000
rect 16200 -8600 18800 -8500
rect 16200 -8900 16300 -8600
rect 18700 -8900 18800 -8600
rect 16200 -9000 18800 -8900
rect 19200 -9200 19600 -300
rect 4900 -9400 19600 -9200
rect 19900 -9400 20000 -100
rect 4500 -9600 20000 -9400
rect 4500 -9900 5100 -9600
rect 19400 -9900 20000 -9600
rect 4500 -10000 20000 -9900
rect -3000 -16500 -2500 -16400
rect 4500 -10600 8500 -10500
rect 4500 -10900 5000 -10600
rect 8000 -10900 8500 -10600
rect 4500 -11000 8500 -10900
rect 4500 -11100 5000 -11000
rect 4500 -15900 4600 -11100
rect 4900 -15900 5000 -11100
rect 8000 -11100 8500 -11000
rect 4500 -16000 5000 -15900
rect 5200 -16000 5700 -12000
rect 8000 -15900 8100 -11100
rect 8400 -15900 8500 -11100
rect 8000 -16000 8500 -15900
rect 4500 -16100 8500 -16000
rect 4500 -16400 5000 -16100
rect 8000 -16400 8500 -16100
rect 4500 -16500 8500 -16400
rect 11500 -10600 20000 -10500
rect 11500 -10900 12100 -10600
rect 19400 -10900 20000 -10600
rect 11500 -11000 20000 -10900
rect 11500 -11100 12000 -11000
rect 11500 -15900 11600 -11100
rect 11900 -15900 12000 -11100
rect 19500 -11100 20000 -11000
rect 11500 -16000 12000 -15900
rect 13900 -16000 14400 -12500
rect 17000 -16000 17500 -12500
rect 19500 -15900 19600 -11100
rect 19900 -15900 20000 -11100
rect 19500 -16000 20000 -15900
rect 11500 -16100 20000 -16000
rect 11500 -16400 12100 -16100
rect 19400 -16400 20000 -16100
rect 11500 -16500 20000 -16400
rect -12000 -16600 -2500 -16500
rect -12000 -16900 -11400 -16600
rect -3100 -16900 -2500 -16600
rect -12000 -17100 -2500 -16900
rect -12000 -17400 -11900 -17100
rect -11600 -17400 -11400 -17100
rect -11100 -17400 -10900 -17100
rect -10600 -17400 -10400 -17100
rect -10100 -17400 -9900 -17100
rect -9600 -17400 -9400 -17100
rect -9100 -17400 -8900 -17100
rect -8600 -17400 -8400 -17100
rect -8100 -17400 -7900 -17100
rect -7600 -17400 -7400 -17100
rect -7100 -17400 -6900 -17100
rect -6600 -17400 -6400 -17100
rect -6100 -17400 -5900 -17100
rect -5600 -17400 -5400 -17100
rect -5100 -17400 -4900 -17100
rect -4600 -17400 -4400 -17100
rect -4100 -17400 -3900 -17100
rect -3600 -17400 -3400 -17100
rect -3100 -17400 -2900 -17100
rect -2600 -17400 -2500 -17100
rect -12000 -17600 -2500 -17400
rect -12000 -17900 -11900 -17600
rect -11600 -17900 -11400 -17600
rect -11100 -17900 -10900 -17600
rect -10600 -17900 -10400 -17600
rect -10100 -17900 -9900 -17600
rect -9600 -17900 -9400 -17600
rect -9100 -17900 -8900 -17600
rect -8600 -17900 -8400 -17600
rect -8100 -17900 -7900 -17600
rect -7600 -17900 -7400 -17600
rect -7100 -17900 -6900 -17600
rect -6600 -17900 -6400 -17600
rect -6100 -17900 -5900 -17600
rect -5600 -17900 -5400 -17600
rect -5100 -17900 -4900 -17600
rect -4600 -17900 -4400 -17600
rect -4100 -17900 -3900 -17600
rect -3600 -17900 -3400 -17600
rect -3100 -17900 -2900 -17600
rect -2600 -17900 -2500 -17600
rect -12000 -18100 -2500 -17900
rect -12000 -18400 -11900 -18100
rect -11600 -18400 -11400 -18100
rect -11100 -18400 -10900 -18100
rect -10600 -18400 -10400 -18100
rect -10100 -18400 -9900 -18100
rect -9600 -18400 -9400 -18100
rect -9100 -18400 -8900 -18100
rect -8600 -18400 -8400 -18100
rect -8100 -18400 -7900 -18100
rect -7600 -18400 -7400 -18100
rect -7100 -18400 -6900 -18100
rect -6600 -18400 -6400 -18100
rect -6100 -18400 -5900 -18100
rect -5600 -18400 -5400 -18100
rect -5100 -18400 -4900 -18100
rect -4600 -18400 -4400 -18100
rect -4100 -18400 -3900 -18100
rect -3600 -18400 -3400 -18100
rect -3100 -18400 -2900 -18100
rect -2600 -18400 -2500 -18100
rect -12000 -18600 -2500 -18400
rect -12000 -18900 -11900 -18600
rect -11600 -18900 -11400 -18600
rect -11100 -18900 -10900 -18600
rect -10600 -18900 -10400 -18600
rect -10100 -18900 -9900 -18600
rect -9600 -18900 -9400 -18600
rect -9100 -18900 -8900 -18600
rect -8600 -18900 -8400 -18600
rect -8100 -18900 -7900 -18600
rect -7600 -18900 -7400 -18600
rect -7100 -18900 -6900 -18600
rect -6600 -18900 -6400 -18600
rect -6100 -18900 -5900 -18600
rect -5600 -18900 -5400 -18600
rect -5100 -18900 -4900 -18600
rect -4600 -18900 -4400 -18600
rect -4100 -18900 -3900 -18600
rect -3600 -18900 -3400 -18600
rect -3100 -18900 -2900 -18600
rect -2600 -18900 -2500 -18600
rect -12000 -19100 -2500 -18900
rect -12000 -19400 -11900 -19100
rect -11600 -19400 -11400 -19100
rect -11100 -19400 -10900 -19100
rect -10600 -19400 -10400 -19100
rect -10100 -19400 -9900 -19100
rect -9600 -19400 -9400 -19100
rect -9100 -19400 -8900 -19100
rect -8600 -19400 -8400 -19100
rect -8100 -19400 -7900 -19100
rect -7600 -19400 -7400 -19100
rect -7100 -19400 -6900 -19100
rect -6600 -19400 -6400 -19100
rect -6100 -19400 -5900 -19100
rect -5600 -19400 -5400 -19100
rect -5100 -19400 -4900 -19100
rect -4600 -19400 -4400 -19100
rect -4100 -19400 -3900 -19100
rect -3600 -19400 -3400 -19100
rect -3100 -19400 -2900 -19100
rect -2600 -19400 -2500 -19100
rect -12000 -19600 -2500 -19400
rect -12000 -19900 -11900 -19600
rect -11600 -19900 -11400 -19600
rect -11100 -19900 -10900 -19600
rect -10600 -19900 -10400 -19600
rect -10100 -19900 -9900 -19600
rect -9600 -19900 -9400 -19600
rect -9100 -19900 -8900 -19600
rect -8600 -19900 -8400 -19600
rect -8100 -19900 -7900 -19600
rect -7600 -19900 -7400 -19600
rect -7100 -19900 -6900 -19600
rect -6600 -19900 -6400 -19600
rect -6100 -19900 -5900 -19600
rect -5600 -19900 -5400 -19600
rect -5100 -19900 -4900 -19600
rect -4600 -19900 -4400 -19600
rect -4100 -19900 -3900 -19600
rect -3600 -19900 -3400 -19600
rect -3100 -19900 -2900 -19600
rect -2600 -19900 -2500 -19600
rect -12000 -20100 -2500 -19900
rect -12000 -20400 -11900 -20100
rect -11600 -20400 -11400 -20100
rect -11100 -20400 -10900 -20100
rect -10600 -20400 -10400 -20100
rect -10100 -20400 -9900 -20100
rect -9600 -20400 -9400 -20100
rect -9100 -20400 -8900 -20100
rect -8600 -20400 -8400 -20100
rect -8100 -20400 -7900 -20100
rect -7600 -20400 -7400 -20100
rect -7100 -20400 -6900 -20100
rect -6600 -20400 -6400 -20100
rect -6100 -20400 -5900 -20100
rect -5600 -20400 -5400 -20100
rect -5100 -20400 -4900 -20100
rect -4600 -20400 -4400 -20100
rect -4100 -20400 -3900 -20100
rect -3600 -20400 -3400 -20100
rect -3100 -20400 -2900 -20100
rect -2600 -20400 -2500 -20100
rect -12000 -20500 -2500 -20400
rect 20500 -26400 20600 6400
rect 20900 -26400 21000 6400
rect 20500 -26500 21000 -26400
rect 23100 -26500 23600 6500
rect 26200 -26500 26700 6500
rect 29000 6400 29500 6500
rect 29000 -26400 29100 6400
rect 29400 -26400 29500 6400
rect 29000 -26500 29500 -26400
rect 20500 -26600 29500 -26500
rect 20500 -26900 21100 -26600
rect 28900 -26900 29500 -26600
rect 20500 -27000 29500 -26900
<< viali >>
rect -11900 10100 -11600 10400
rect -11900 9600 -11600 9900
rect -11900 9100 -11600 9400
rect -11900 8600 -11600 8900
rect -11900 8100 -11600 8400
rect -11900 7600 -11600 7900
rect -11900 7100 -11600 7400
rect 12100 -900 12400 -600
rect 12100 -1400 12400 -1100
rect 12100 -1900 12400 -1600
rect 12100 -2400 12400 -2100
rect 12100 -2900 12400 -2600
rect 12100 -3400 12400 -3100
rect 12100 -6400 12400 -6100
rect 12100 -6900 12400 -6600
rect 12100 -7400 12400 -7100
rect 12100 -7900 12400 -7600
rect 12100 -8400 12400 -8100
rect 12100 -8900 12400 -8600
rect -11900 -17400 -11600 -17100
rect -11400 -17400 -11100 -17100
rect -10900 -17400 -10600 -17100
rect -10400 -17400 -10100 -17100
rect -9900 -17400 -9600 -17100
rect -9400 -17400 -9100 -17100
rect -8900 -17400 -8600 -17100
rect -8400 -17400 -8100 -17100
rect -7900 -17400 -7600 -17100
rect -7400 -17400 -7100 -17100
rect -6900 -17400 -6600 -17100
rect -6400 -17400 -6100 -17100
rect -5900 -17400 -5600 -17100
rect -5400 -17400 -5100 -17100
rect -4900 -17400 -4600 -17100
rect -4400 -17400 -4100 -17100
rect -3900 -17400 -3600 -17100
rect -3400 -17400 -3100 -17100
rect -2900 -17400 -2600 -17100
rect -11900 -17900 -11600 -17600
rect -11400 -17900 -11100 -17600
rect -10900 -17900 -10600 -17600
rect -10400 -17900 -10100 -17600
rect -9900 -17900 -9600 -17600
rect -9400 -17900 -9100 -17600
rect -8900 -17900 -8600 -17600
rect -8400 -17900 -8100 -17600
rect -7900 -17900 -7600 -17600
rect -7400 -17900 -7100 -17600
rect -6900 -17900 -6600 -17600
rect -6400 -17900 -6100 -17600
rect -5900 -17900 -5600 -17600
rect -5400 -17900 -5100 -17600
rect -4900 -17900 -4600 -17600
rect -4400 -17900 -4100 -17600
rect -3900 -17900 -3600 -17600
rect -3400 -17900 -3100 -17600
rect -2900 -17900 -2600 -17600
rect -11900 -18400 -11600 -18100
rect -11400 -18400 -11100 -18100
rect -10900 -18400 -10600 -18100
rect -10400 -18400 -10100 -18100
rect -9900 -18400 -9600 -18100
rect -9400 -18400 -9100 -18100
rect -8900 -18400 -8600 -18100
rect -8400 -18400 -8100 -18100
rect -7900 -18400 -7600 -18100
rect -7400 -18400 -7100 -18100
rect -6900 -18400 -6600 -18100
rect -6400 -18400 -6100 -18100
rect -5900 -18400 -5600 -18100
rect -5400 -18400 -5100 -18100
rect -4900 -18400 -4600 -18100
rect -4400 -18400 -4100 -18100
rect -3900 -18400 -3600 -18100
rect -3400 -18400 -3100 -18100
rect -2900 -18400 -2600 -18100
rect -11900 -18900 -11600 -18600
rect -11400 -18900 -11100 -18600
rect -10900 -18900 -10600 -18600
rect -10400 -18900 -10100 -18600
rect -9900 -18900 -9600 -18600
rect -9400 -18900 -9100 -18600
rect -8900 -18900 -8600 -18600
rect -8400 -18900 -8100 -18600
rect -7900 -18900 -7600 -18600
rect -7400 -18900 -7100 -18600
rect -6900 -18900 -6600 -18600
rect -6400 -18900 -6100 -18600
rect -5900 -18900 -5600 -18600
rect -5400 -18900 -5100 -18600
rect -4900 -18900 -4600 -18600
rect -4400 -18900 -4100 -18600
rect -3900 -18900 -3600 -18600
rect -3400 -18900 -3100 -18600
rect -2900 -18900 -2600 -18600
rect -11900 -19400 -11600 -19100
rect -11400 -19400 -11100 -19100
rect -10900 -19400 -10600 -19100
rect -10400 -19400 -10100 -19100
rect -9900 -19400 -9600 -19100
rect -9400 -19400 -9100 -19100
rect -8900 -19400 -8600 -19100
rect -8400 -19400 -8100 -19100
rect -7900 -19400 -7600 -19100
rect -7400 -19400 -7100 -19100
rect -6900 -19400 -6600 -19100
rect -6400 -19400 -6100 -19100
rect -5900 -19400 -5600 -19100
rect -5400 -19400 -5100 -19100
rect -4900 -19400 -4600 -19100
rect -4400 -19400 -4100 -19100
rect -3900 -19400 -3600 -19100
rect -3400 -19400 -3100 -19100
rect -2900 -19400 -2600 -19100
rect -11900 -19900 -11600 -19600
rect -11400 -19900 -11100 -19600
rect -10900 -19900 -10600 -19600
rect -10400 -19900 -10100 -19600
rect -9900 -19900 -9600 -19600
rect -9400 -19900 -9100 -19600
rect -8900 -19900 -8600 -19600
rect -8400 -19900 -8100 -19600
rect -7900 -19900 -7600 -19600
rect -7400 -19900 -7100 -19600
rect -6900 -19900 -6600 -19600
rect -6400 -19900 -6100 -19600
rect -5900 -19900 -5600 -19600
rect -5400 -19900 -5100 -19600
rect -4900 -19900 -4600 -19600
rect -4400 -19900 -4100 -19600
rect -3900 -19900 -3600 -19600
rect -3400 -19900 -3100 -19600
rect -2900 -19900 -2600 -19600
rect -11900 -20400 -11600 -20100
rect -11400 -20400 -11100 -20100
rect -10900 -20400 -10600 -20100
rect -10400 -20400 -10100 -20100
rect -9900 -20400 -9600 -20100
rect -9400 -20400 -9100 -20100
rect -8900 -20400 -8600 -20100
rect -8400 -20400 -8100 -20100
rect -7900 -20400 -7600 -20100
rect -7400 -20400 -7100 -20100
rect -6900 -20400 -6600 -20100
rect -6400 -20400 -6100 -20100
rect -5900 -20400 -5600 -20100
rect -5400 -20400 -5100 -20100
rect -4900 -20400 -4600 -20100
rect -4400 -20400 -4100 -20100
rect -3900 -20400 -3600 -20100
rect -3400 -20400 -3100 -20100
rect -2900 -20400 -2600 -20100
<< metal1 >>
rect -12000 10400 -2500 10500
rect -12000 10100 -11900 10400
rect -11600 10100 -2500 10400
rect -12000 9900 -2500 10100
rect -12000 9600 -11900 9900
rect -11600 9600 -2500 9900
rect -12000 9400 -2500 9600
rect -12000 9100 -11900 9400
rect -11600 9100 -2500 9400
rect -12000 8900 -2500 9100
rect -12000 8600 -11900 8900
rect -11600 8600 -2500 8900
rect -12000 8400 -2500 8600
rect -12000 8100 -11900 8400
rect -11600 8100 -2500 8400
rect -12000 7900 -2500 8100
rect -12000 7600 -11900 7900
rect -11600 7600 -2500 7900
rect -12000 7400 -2500 7600
rect -12000 7100 -11900 7400
rect -11600 7100 -2500 7400
rect -12000 7000 -2500 7100
rect -10900 4400 -10400 4500
rect -10900 4100 -10800 4400
rect -10500 4100 -10400 4400
rect -10900 3900 -10400 4100
rect -10900 3600 -10800 3900
rect -10500 3600 -10400 3900
rect -10900 3500 -10400 3600
rect -7800 4400 -7300 4500
rect -7800 4100 -7700 4400
rect -7400 4100 -7300 4400
rect -7800 3900 -7300 4100
rect -7800 3600 -7700 3900
rect -7400 3600 -7300 3900
rect -7800 3500 -7300 3600
rect -4700 4400 -4200 4500
rect -4700 4100 -4600 4400
rect -4300 4100 -4200 4400
rect -4700 3900 -4200 4100
rect -4700 3600 -4600 3900
rect -4300 3600 -4200 3900
rect -4700 3500 -4200 3600
rect -3900 2300 -3400 5200
rect -900 2300 -400 5200
rect 2200 2300 2700 5200
rect -11000 1800 2700 2300
rect 6000 2500 6500 5500
rect 8900 4400 9500 4500
rect 8900 4100 9000 4400
rect 9300 4100 9500 4400
rect 8900 3900 9500 4100
rect 8900 3600 9000 3900
rect 9300 3600 9500 3900
rect 8900 3500 9500 3600
rect 12000 2500 12500 5500
rect 15100 4400 15700 4500
rect 15100 4100 15300 4400
rect 15600 4100 15700 4400
rect 15100 3900 15700 4100
rect 15100 3600 15300 3900
rect 15600 3600 15700 3900
rect 15100 3500 15700 3600
rect 18000 2500 18500 5500
rect 6000 2000 18500 2500
rect 20000 5000 28000 6000
rect 20000 4400 21000 5000
rect 20000 4100 20100 4400
rect 20400 4100 20600 4400
rect 20900 4100 21000 4400
rect 20000 3900 21000 4100
rect 20000 3600 20100 3900
rect 20400 3600 20600 3900
rect 20900 3600 21000 3900
rect -9700 -1700 -9200 1800
rect -10200 -2000 -9200 -1700
rect -9700 -2200 -9200 -2000
rect -10900 -4500 -10400 -2200
rect -9900 -3100 -9200 -2200
rect -9700 -3300 -9200 -3100
rect -10200 -3600 -9200 -3300
rect -6700 1400 -6200 1500
rect -6700 1100 -6600 1400
rect -6300 1100 -6200 1400
rect -6700 900 -6200 1100
rect -6700 600 -6600 900
rect -6300 600 -6200 900
rect -6700 -4500 -6200 600
rect -10900 -4700 -6200 -4500
rect -4500 -4600 -3300 -1200
rect -1900 -4600 -1400 1800
rect 20000 400 21000 3600
rect 21700 2000 22200 3000
rect 24600 2000 25100 3000
rect 27700 2000 28200 3000
rect 20000 100 20100 400
rect 20400 100 20600 400
rect 20900 100 21000 400
rect 20000 0 21000 100
rect 20000 -100 28000 0
rect 20000 -400 20100 -100
rect 20400 -400 20600 -100
rect 20900 -400 28000 -100
rect 12050 -600 12450 -500
rect 12050 -900 12100 -600
rect 12400 -900 12450 -600
rect 12050 -1100 12450 -900
rect 20000 -1000 28000 -400
rect 10200 -1600 10700 -1300
rect 12000 -1400 12100 -1100
rect 12400 -1400 12500 -1100
rect 12000 -1600 12500 -1400
rect 13700 -1600 14200 -1300
rect 12050 -1900 12100 -1600
rect 12400 -1900 12450 -1600
rect 7200 -3000 8000 -1900
rect 8500 -2100 9000 -2000
rect 8500 -2400 8600 -2100
rect 8900 -2400 9000 -2100
rect 8500 -2500 9000 -2400
rect 8500 -2800 8600 -2500
rect 8900 -2800 9000 -2500
rect 8500 -2900 9000 -2800
rect 8500 -3200 8600 -2900
rect 8900 -3200 9000 -2900
rect 9400 -3000 10200 -1900
rect 12050 -2100 12450 -1900
rect 12050 -2400 12100 -2100
rect 12400 -2400 12450 -2100
rect 12050 -2600 12450 -2400
rect 12050 -2900 12100 -2600
rect 12400 -2900 12450 -2600
rect 12050 -3050 12450 -2900
rect 14100 -3000 14900 -1900
rect 16500 -3000 17300 -1900
rect 6700 -4000 7200 -3200
rect 8500 -3300 9000 -3200
rect 8500 -3600 8600 -3300
rect 8900 -3600 9000 -3300
rect 11100 -3100 13400 -3050
rect 11100 -3400 11150 -3100
rect 11450 -3400 12100 -3100
rect 12400 -3400 13050 -3100
rect 13350 -3400 13400 -3100
rect 11100 -3450 13400 -3400
rect 8500 -3700 9000 -3600
rect 8500 -4000 8600 -3700
rect 8900 -4000 9000 -3700
rect 12050 -3800 12450 -3450
rect 17200 -4000 17700 -3200
rect 500 -4100 19500 -4000
rect 500 -4400 8600 -4100
rect 8900 -4400 19500 -4100
rect 500 -4500 19500 -4400
rect -10900 -5000 -5000 -4700
rect -6200 -6000 -5000 -5000
rect -11000 -10000 -9000 -8500
rect -4500 -8900 -3700 -4600
rect -3200 -6000 -2000 -4700
rect -4100 -9100 -3600 -8900
rect -5500 -12000 -3500 -10500
rect -11000 -13500 -9000 -12000
rect -5500 -15000 -3500 -13500
rect -12000 -17100 -2500 -17000
rect -12000 -17400 -11900 -17100
rect -11600 -17400 -11400 -17100
rect -11100 -17400 -10900 -17100
rect -10600 -17400 -10400 -17100
rect -10100 -17400 -9900 -17100
rect -9600 -17400 -9400 -17100
rect -9100 -17400 -8900 -17100
rect -8600 -17400 -8400 -17100
rect -8100 -17400 -7900 -17100
rect -7600 -17400 -7400 -17100
rect -7100 -17400 -6900 -17100
rect -6600 -17400 -6400 -17100
rect -6100 -17400 -5900 -17100
rect -5600 -17400 -5400 -17100
rect -5100 -17400 -4900 -17100
rect -4600 -17400 -4400 -17100
rect -4100 -17400 -3900 -17100
rect -3600 -17400 -3400 -17100
rect -3100 -17400 -2900 -17100
rect -2600 -17400 -2500 -17100
rect -12000 -17600 -2500 -17400
rect -12000 -17900 -11900 -17600
rect -11600 -17900 -11400 -17600
rect -11100 -17900 -10900 -17600
rect -10600 -17900 -10400 -17600
rect -10100 -17900 -9900 -17600
rect -9600 -17900 -9400 -17600
rect -9100 -17900 -8900 -17600
rect -8600 -17900 -8400 -17600
rect -8100 -17900 -7900 -17600
rect -7600 -17900 -7400 -17600
rect -7100 -17900 -6900 -17600
rect -6600 -17900 -6400 -17600
rect -6100 -17900 -5900 -17600
rect -5600 -17900 -5400 -17600
rect -5100 -17900 -4900 -17600
rect -4600 -17900 -4400 -17600
rect -4100 -17900 -3900 -17600
rect -3600 -17900 -3400 -17600
rect -3100 -17900 -2900 -17600
rect -2600 -17900 -2500 -17600
rect -12000 -18100 -2500 -17900
rect -12000 -18400 -11900 -18100
rect -11600 -18400 -11400 -18100
rect -11100 -18400 -10900 -18100
rect -10600 -18400 -10400 -18100
rect -10100 -18400 -9900 -18100
rect -9600 -18400 -9400 -18100
rect -9100 -18400 -8900 -18100
rect -8600 -18400 -8400 -18100
rect -8100 -18400 -7900 -18100
rect -7600 -18400 -7400 -18100
rect -7100 -18400 -6900 -18100
rect -6600 -18400 -6400 -18100
rect -6100 -18400 -5900 -18100
rect -5600 -18400 -5400 -18100
rect -5100 -18400 -4900 -18100
rect -4600 -18400 -4400 -18100
rect -4100 -18400 -3900 -18100
rect -3600 -18400 -3400 -18100
rect -3100 -18400 -2900 -18100
rect -2600 -18400 -2500 -18100
rect -12000 -18600 -2500 -18400
rect -12000 -18900 -11900 -18600
rect -11600 -18900 -11400 -18600
rect -11100 -18900 -10900 -18600
rect -10600 -18900 -10400 -18600
rect -10100 -18900 -9900 -18600
rect -9600 -18900 -9400 -18600
rect -9100 -18900 -8900 -18600
rect -8600 -18900 -8400 -18600
rect -8100 -18900 -7900 -18600
rect -7600 -18900 -7400 -18600
rect -7100 -18900 -6900 -18600
rect -6600 -18900 -6400 -18600
rect -6100 -18900 -5900 -18600
rect -5600 -18900 -5400 -18600
rect -5100 -18900 -4900 -18600
rect -4600 -18900 -4400 -18600
rect -4100 -18900 -3900 -18600
rect -3600 -18900 -3400 -18600
rect -3100 -18900 -2900 -18600
rect -2600 -18900 -2500 -18600
rect -12000 -19100 -2500 -18900
rect -12000 -19400 -11900 -19100
rect -11600 -19400 -11400 -19100
rect -11100 -19400 -10900 -19100
rect -10600 -19400 -10400 -19100
rect -10100 -19400 -9900 -19100
rect -9600 -19400 -9400 -19100
rect -9100 -19400 -8900 -19100
rect -8600 -19400 -8400 -19100
rect -8100 -19400 -7900 -19100
rect -7600 -19400 -7400 -19100
rect -7100 -19400 -6900 -19100
rect -6600 -19400 -6400 -19100
rect -6100 -19400 -5900 -19100
rect -5600 -19400 -5400 -19100
rect -5100 -19400 -4900 -19100
rect -4600 -19400 -4400 -19100
rect -4100 -19400 -3900 -19100
rect -3600 -19400 -3400 -19100
rect -3100 -19400 -2900 -19100
rect -2600 -19400 -2500 -19100
rect -12000 -19600 -2500 -19400
rect -12000 -19900 -11900 -19600
rect -11600 -19900 -11400 -19600
rect -11100 -19900 -10900 -19600
rect -10600 -19900 -10400 -19600
rect -10100 -19900 -9900 -19600
rect -9600 -19900 -9400 -19600
rect -9100 -19900 -8900 -19600
rect -8600 -19900 -8400 -19600
rect -8100 -19900 -7900 -19600
rect -7600 -19900 -7400 -19600
rect -7100 -19900 -6900 -19600
rect -6600 -19900 -6400 -19600
rect -6100 -19900 -5900 -19600
rect -5600 -19900 -5400 -19600
rect -5100 -19900 -4900 -19600
rect -4600 -19900 -4400 -19600
rect -4100 -19900 -3900 -19600
rect -3600 -19900 -3400 -19600
rect -3100 -19900 -2900 -19600
rect -2600 -19900 -2500 -19600
rect -12000 -20100 -2500 -19900
rect -12000 -20400 -11900 -20100
rect -11600 -20400 -11400 -20100
rect -11100 -20400 -10900 -20100
rect -10600 -20400 -10400 -20100
rect -10100 -20400 -9900 -20100
rect -9600 -20400 -9400 -20100
rect -9100 -20400 -8900 -20100
rect -8600 -20400 -8400 -20100
rect -8100 -20400 -7900 -20100
rect -7600 -20400 -7400 -20100
rect -7100 -20400 -6900 -20100
rect -6600 -20400 -6400 -20100
rect -6100 -20400 -5900 -20100
rect -5600 -20400 -5400 -20100
rect -5100 -20400 -4900 -20100
rect -4600 -20400 -4400 -20100
rect -4100 -20400 -3900 -20100
rect -3600 -20400 -3400 -20100
rect -3100 -20400 -2900 -20100
rect -2600 -20400 -2500 -20100
rect -12000 -20500 -2500 -20400
rect 500 -21900 1000 -4500
rect 15500 -5000 15600 -4900
rect 2000 -5200 15600 -5000
rect 15900 -5000 16000 -4900
rect 15900 -5200 19500 -5000
rect 2000 -5300 19500 -5200
rect 2000 -5500 15600 -5300
rect 2000 -21900 2500 -5500
rect 6700 -6200 7200 -5500
rect 15500 -5600 15600 -5500
rect 15900 -5500 19500 -5300
rect 15900 -5600 16000 -5500
rect 15500 -5700 16000 -5600
rect 12050 -5950 12450 -5700
rect 11100 -6000 13400 -5950
rect 11100 -6300 11150 -6000
rect 11450 -6100 13050 -6000
rect 11450 -6300 12100 -6100
rect 11100 -6350 12100 -6300
rect 12050 -6400 12100 -6350
rect 12400 -6300 13050 -6100
rect 13350 -6300 13400 -6000
rect 12400 -6350 13400 -6300
rect 15500 -6000 15600 -5700
rect 15900 -6000 16000 -5700
rect 15500 -6100 16000 -6000
rect 12400 -6400 12450 -6350
rect 15500 -6400 15600 -6100
rect 15900 -6400 16000 -6100
rect 17200 -6200 17700 -5500
rect 6000 -7500 6800 -6400
rect 9500 -7500 10300 -6400
rect 12050 -6600 12450 -6400
rect 12050 -6900 12100 -6600
rect 12400 -6900 12450 -6600
rect 12050 -7100 12450 -6900
rect 12050 -7400 12100 -7100
rect 12400 -7400 12450 -7100
rect 12050 -7600 12450 -7400
rect 14100 -7500 14900 -6400
rect 15500 -6500 16000 -6400
rect 15500 -6800 15600 -6500
rect 15900 -6800 16000 -6500
rect 15500 -6900 16000 -6800
rect 15500 -7200 15600 -6900
rect 15900 -7200 16000 -6900
rect 15500 -7300 16000 -7200
rect 17600 -7500 18400 -6400
rect 20000 -6500 21000 -1000
rect 21700 -4400 22200 -3400
rect 24700 -4400 25200 -3400
rect 27700 -4400 28200 -3400
rect 20000 -7500 28000 -6500
rect 12050 -7700 12100 -7600
rect 10200 -8000 10700 -7700
rect 12000 -7900 12100 -7700
rect 12400 -7700 12450 -7600
rect 12400 -7900 12500 -7700
rect 12000 -8100 12500 -7900
rect 13700 -8000 14200 -7700
rect 12000 -8200 12100 -8100
rect 12050 -8400 12100 -8200
rect 12400 -8200 12500 -8100
rect 12400 -8400 12450 -8200
rect 12050 -8500 12450 -8400
rect 12000 -8600 12500 -8500
rect 12000 -8900 12100 -8600
rect 12400 -8900 12500 -8600
rect 12000 -10000 12500 -8900
rect 9700 -10400 12500 -10000
rect 20000 -9100 21000 -7500
rect 20000 -9400 20100 -9100
rect 20400 -9400 20600 -9100
rect 20900 -9400 21000 -9100
rect 20000 -9600 21000 -9400
rect 20000 -9900 20100 -9600
rect 20400 -9900 20600 -9600
rect 20900 -9900 21000 -9600
rect 7100 -16000 7600 -12000
rect 9700 -16000 10200 -10400
rect 20000 -13000 21000 -9900
rect 21700 -10800 22200 -9800
rect 24700 -10800 25200 -9800
rect 27700 -10800 28200 -9800
rect 12500 -14500 13000 -13500
rect 15500 -14500 16000 -13500
rect 18600 -14500 19100 -13500
rect 20000 -14000 28000 -13000
rect 7100 -16500 10200 -16000
rect 20000 -19000 21000 -14000
rect 21700 -17200 22200 -16200
rect 24600 -17200 25100 -16200
rect 27700 -17200 28200 -16200
rect 20000 -20000 28000 -19000
rect 200 -22900 1200 -21900
rect 1800 -22900 2800 -21900
rect 21700 -23500 22200 -22500
rect 24600 -23500 25100 -22500
rect 27700 -23500 28200 -22500
rect 18500 -25600 19500 -25500
rect 18500 -25900 18600 -25600
rect 18900 -25900 19100 -25600
rect 19400 -25900 19500 -25600
rect 18500 -26100 19500 -25900
rect 18500 -26400 18600 -26100
rect 18900 -26400 19100 -26100
rect 19400 -26400 19500 -26100
rect 18500 -26500 19500 -26400
<< via1 >>
rect -10800 4100 -10500 4400
rect -10800 3600 -10500 3900
rect -7700 4100 -7400 4400
rect -7700 3600 -7400 3900
rect -4600 4100 -4300 4400
rect -4600 3600 -4300 3900
rect 9000 4100 9300 4400
rect 9000 3600 9300 3900
rect 15300 4100 15600 4400
rect 15300 3600 15600 3900
rect 20100 4100 20400 4400
rect 20600 4100 20900 4400
rect 20100 3600 20400 3900
rect 20600 3600 20900 3900
rect -6600 1100 -6300 1400
rect -6600 600 -6300 900
rect 20100 100 20400 400
rect 20600 100 20900 400
rect 20100 -400 20400 -100
rect 20600 -400 20900 -100
rect 8600 -2400 8900 -2100
rect 8600 -2800 8900 -2500
rect 8600 -3200 8900 -2900
rect 8600 -3600 8900 -3300
rect 11150 -3400 11450 -3100
rect 13050 -3400 13350 -3100
rect 8600 -4000 8900 -3700
rect 8600 -4400 8900 -4100
rect 15600 -5200 15900 -4900
rect 15600 -5600 15900 -5300
rect 11150 -6300 11450 -6000
rect 13050 -6300 13350 -6000
rect 15600 -6000 15900 -5700
rect 15600 -6400 15900 -6100
rect 15600 -6800 15900 -6500
rect 15600 -7200 15900 -6900
rect 20100 -9400 20400 -9100
rect 20600 -9400 20900 -9100
rect 20100 -9900 20400 -9600
rect 20600 -9900 20900 -9600
rect 18600 -25900 18900 -25600
rect 19100 -25900 19400 -25600
rect 18600 -26400 18900 -26100
rect 19100 -26400 19400 -26100
<< metal2 >>
rect -11500 4400 -4000 4500
rect -11500 4100 -10800 4400
rect -10500 4100 -7700 4400
rect -7400 4100 -4600 4400
rect -4300 4100 -4000 4400
rect -11500 3900 -4000 4100
rect -11500 3600 -10800 3900
rect -10500 3600 -7700 3900
rect -7400 3600 -4600 3900
rect -4300 3600 -4000 3900
rect -11500 3500 -4000 3600
rect 5500 4400 21000 4500
rect 5500 4100 9000 4400
rect 9300 4100 15300 4400
rect 15600 4100 20100 4400
rect 20400 4100 20600 4400
rect 20900 4100 21000 4400
rect 5500 3900 21000 4100
rect 5500 3600 9000 3900
rect 9300 3600 15300 3900
rect 15600 3600 20100 3900
rect 20400 3600 20600 3900
rect 20900 3600 21000 3900
rect 5500 3500 21000 3600
rect -8000 1500 -7200 3500
rect 21700 2000 29500 3000
rect -10500 1400 2500 1500
rect -10500 1100 -6600 1400
rect -6300 1100 2500 1400
rect -10500 900 2500 1100
rect 5000 1000 19500 2000
rect -10500 600 -6600 900
rect -6300 600 2500 900
rect -10500 500 2500 600
rect 5500 400 21000 500
rect 5500 100 20100 400
rect 20400 100 20600 400
rect 20900 100 21000 400
rect 5500 -100 21000 100
rect 5500 -400 20100 -100
rect 20400 -400 20600 -100
rect 20900 -400 21000 -100
rect 5500 -500 21000 -400
rect -6500 -6000 0 -5000
rect -1000 -10500 0 -6000
rect 6000 -6400 6500 -1000
rect 9300 -1900 9800 -500
rect 10000 -1600 16000 -1100
rect 7200 -3000 8000 -1900
rect 8500 -2100 9000 -2000
rect 8500 -2400 8600 -2100
rect 8900 -2400 9000 -2100
rect 8500 -2500 9000 -2400
rect 8500 -2800 8600 -2500
rect 8900 -2800 9000 -2500
rect 8500 -2900 9000 -2800
rect 8500 -3200 8600 -2900
rect 8900 -3200 9000 -2900
rect 8500 -3300 9000 -3200
rect 8500 -3600 8600 -3300
rect 8900 -3600 9000 -3300
rect 8500 -3700 9000 -3600
rect 8500 -4000 8600 -3700
rect 8900 -4000 9000 -3700
rect 9300 -2200 10200 -1900
rect 14100 -2200 14900 -1900
rect 9300 -2700 14900 -2200
rect 9300 -3000 10200 -2700
rect 14100 -3000 14900 -2700
rect 9300 -4000 9800 -3000
rect 11100 -3100 11500 -3050
rect 11100 -3400 11150 -3100
rect 11450 -3400 11500 -3100
rect 11100 -3450 11500 -3400
rect 13000 -3100 13400 -3050
rect 13000 -3400 13050 -3100
rect 13350 -3400 13400 -3100
rect 13000 -3450 13400 -3400
rect 8500 -4100 9000 -4000
rect 8500 -4400 8600 -4100
rect 8900 -4400 9000 -4100
rect 6000 -7500 6800 -6400
rect 6000 -9000 6500 -7500
rect 8500 -7700 9000 -4400
rect 15500 -4900 16000 -1600
rect 16500 -3000 17300 -1900
rect 15500 -5200 15600 -4900
rect 15900 -5200 16000 -4900
rect 15500 -5300 16000 -5200
rect 15500 -5600 15600 -5300
rect 15900 -5600 16000 -5300
rect 15500 -5700 16000 -5600
rect 11100 -6000 11500 -5950
rect 11100 -6300 11150 -6000
rect 11450 -6300 11500 -6000
rect 11100 -6350 11500 -6300
rect 13000 -6000 13400 -5950
rect 13000 -6300 13050 -6000
rect 13350 -6300 13400 -6000
rect 13000 -6350 13400 -6300
rect 15500 -6000 15600 -5700
rect 15900 -6000 16000 -5700
rect 15500 -6100 16000 -6000
rect 15500 -6400 15600 -6100
rect 15900 -6400 16000 -6100
rect 18000 -6400 18500 -1000
rect 28600 -3400 29500 2000
rect 21700 -4400 29500 -3400
rect 9500 -7500 10300 -6400
rect 14100 -7500 15000 -6400
rect 15500 -6500 16000 -6400
rect 15500 -6800 15600 -6500
rect 15900 -6800 16000 -6500
rect 15500 -6900 16000 -6800
rect 15500 -7200 15600 -6900
rect 15900 -7200 16000 -6900
rect 15500 -7300 16000 -7200
rect 17600 -7500 18500 -6400
rect 8500 -8200 14500 -7700
rect 18000 -9000 18500 -7500
rect 5500 -9100 21000 -9000
rect 5500 -9400 20100 -9100
rect 20400 -9400 20600 -9100
rect 20900 -9400 21000 -9100
rect 5500 -9600 21000 -9400
rect 5500 -9900 20100 -9600
rect 20400 -9900 20600 -9600
rect 20900 -9900 21000 -9600
rect 28600 -9800 29500 -4400
rect 5500 -10000 21000 -9900
rect -1000 -11500 19500 -10500
rect 21700 -10800 29500 -9800
rect 28600 -13500 29500 -10800
rect 12500 -14500 29500 -13500
rect 28600 -16200 29500 -14500
rect 21700 -17200 29500 -16200
rect 28600 -22500 29500 -17200
rect 21700 -23500 29500 -22500
rect 28600 -25500 29500 -23500
rect 18500 -25600 29500 -25500
rect 18500 -25900 18600 -25600
rect 18900 -25900 19100 -25600
rect 19400 -25900 29500 -25600
rect 18500 -26100 29500 -25900
rect 18500 -26400 18600 -26100
rect 18900 -26400 19100 -26100
rect 19400 -26400 29500 -26100
rect 18500 -26500 29500 -26400
<< via2 >>
rect 11150 -3400 11450 -3100
rect 13050 -3400 13350 -3100
rect 11150 -6300 11450 -6000
rect 13050 -6300 13350 -6000
<< metal3 >>
rect 7500 -8000 8000 1500
rect 9500 -8000 10000 1500
rect 11100 -3100 11500 -3050
rect 11100 -3400 11150 -3100
rect 11450 -3400 11500 -3100
rect 11100 -6000 11500 -3400
rect 11100 -6300 11150 -6000
rect 11450 -6300 11500 -6000
rect 11100 -6350 11500 -6300
rect 13000 -3100 13400 -3050
rect 13000 -3400 13050 -3100
rect 13350 -3400 13400 -3100
rect 13000 -6000 13400 -3400
rect 13000 -6300 13050 -6000
rect 13350 -6300 13400 -6000
rect 13000 -6350 13400 -6300
rect 14500 -8000 15000 1500
rect 16500 -8000 17000 1500
<< metal4 >>
rect 20000 7500 48500 8500
rect 30000 -27000 31000 7500
rect 39000 -27500 40000 6500
rect 47500 -27000 48500 7500
rect 57000 -27500 58000 6500
rect 20000 -28500 58000 -27500
use pfet_03v3_SEKV7M  pfet_03v3_SEKV7M_0
timestamp 1771420802
transform 1 0 29350 0 1 27910
box -4590 -16580 4590 16580
use sky130_fd_pr__cap_mim_m3_1_HGK9NV  sky130_fd_pr__cap_mim_m3_1_HGK9NV_0
timestamp 1771414049
transform -1 0 47460 0 -1 -10400
box -17460 -16600 17460 16600
use sky130_fd_pr__nfet_01v8_7PHSG7  sky130_fd_pr__nfet_01v8_7PHSG7_0
timestamp 1771413069
transform 1 0 6940 0 1 -6935
box -440 -1065 440 1065
use sky130_fd_pr__nfet_01v8_7PHSG7  sky130_fd_pr__nfet_01v8_7PHSG7_1
timestamp 1771413069
transform 1 0 13940 0 1 -2435
box -440 -1065 440 1065
use sky130_fd_pr__nfet_01v8_7PHSG7  sky130_fd_pr__nfet_01v8_7PHSG7_2
timestamp 1771413069
transform 1 0 17440 0 1 -2435
box -440 -1065 440 1065
use sky130_fd_pr__nfet_01v8_7PHSG7  sky130_fd_pr__nfet_01v8_7PHSG7_3
timestamp 1771413069
transform 1 0 10440 0 1 -6935
box -440 -1065 440 1065
use sky130_fd_pr__nfet_01v8_7PHSG7  sky130_fd_pr__nfet_01v8_7PHSG7_4
timestamp 1771413069
transform 1 0 10440 0 1 -2435
box -440 -1065 440 1065
use sky130_fd_pr__nfet_01v8_7PHSG7  sky130_fd_pr__nfet_01v8_7PHSG7_5
timestamp 1771413069
transform 1 0 13940 0 1 -6935
box -440 -1065 440 1065
use sky130_fd_pr__nfet_01v8_7PHSG7  sky130_fd_pr__nfet_01v8_7PHSG7_6
timestamp 1771413069
transform 1 0 17440 0 1 -6935
box -440 -1065 440 1065
use sky130_fd_pr__nfet_01v8_K99WZJ  sky130_fd_pr__nfet_01v8_K99WZJ_0
timestamp 1771414049
transform 1 0 -5585 0 1 -3015
box -915 -1985 915 1985
use sky130_fd_pr__pfet_01v8_E2QEAN  sky130_fd_pr__pfet_01v8_E2QEAN_0
timestamp 1771413069
transform 1 0 -7595 0 1 3670
box -3405 -1670 3405 1840
use sky130_fd_pr__res_high_po_1p41_Z9HR6K  sky130_fd_pr__res_high_po_1p41_Z9HR6K_0
timestamp 1771413069
transform 0 1 -7300 -1 0 -10095
box -705 -3700 705 3700
use sky130_fd_pr__res_high_po_1p41_Z9HR6K  sky130_fd_pr__res_high_po_1p41_Z9HR6K_1
timestamp 1771413069
transform 0 1 -7300 -1 0 -11795
box -705 -3700 705 3700
use sky130_fd_pr__res_high_po_1p41_Z9HR6K  sky130_fd_pr__res_high_po_1p41_Z9HR6K_2
timestamp 1771413069
transform 0 1 -7300 -1 0 -13495
box -705 -3700 705 3700
use sky130_fd_pr__res_high_po_1p41_Z9HR6K  sky130_fd_pr__res_high_po_1p41_Z9HR6K_3
timestamp 1771413069
transform 0 1 -7300 -1 0 -15195
box -705 -3700 705 3700
use sky130_fd_pr__nfet_01v8_7PHSG7  XM2
timestamp 1771413069
transform 1 0 6940 0 1 -2435
box -440 -1065 440 1065
use sky130_fd_pr__pfet_01v8_ES843Y  XM4
timestamp 1771413069
transform 1 0 12285 0 1 3870
box -6485 -1670 6485 1840
use sky130_fd_pr__nfet_01v8_K99WZJ  XM5
timestamp 1771414049
transform 1 0 -2585 0 1 -3015
box -915 -1985 915 1985
use sky130_fd_pr__nfet_01v8_68987S  XM7
timestamp 1771413069
transform -1 0 15725 0 -1 -13715
box -3225 -1785 3225 1785
use sky130_fd_pr__pfet_01v8_E2QEAN  XM8
timestamp 1771413069
transform 1 0 -595 0 1 3670
box -3405 -1670 3405 1840
use sky130_fd_pr__nfet_01v8_3RG5EU  XM9
timestamp 1771413069
transform 1 0 6415 0 1 -13515
box -915 -1985 915 1985
use sky130_fd_pr__nfet_01v8_TYFUKG  XM12
timestamp 1771413069
transform 1 0 -10135 0 1 -2635
box -365 -865 365 865
use sky130_fd_pr__res_high_po_1p41_Z9HR6K  XR6
timestamp 1771413069
transform 0 1 -7300 -1 0 -8395
box -705 -3700 705 3700
<< labels >>
flabel metal1 200 -22900 1200 -21900 0 FreeSans 1280 0 0 0 VP
port 2 nsew
flabel metal1 1800 -22900 2800 -21900 0 FreeSans 1280 0 0 0 VN
port 3 nsew
flabel metal1 -8700 7600 -7700 8600 0 FreeSans 1280 0 0 0 VDD
port 0 nsew
flabel metal1 18500 -26500 19500 -25500 0 FreeSans 1280 0 0 0 OUT
port 1 nsew
flabel metal1 -7700 -19000 -6700 -18000 0 FreeSans 1280 0 0 0 VSS
port 4 nsew
<< end >>

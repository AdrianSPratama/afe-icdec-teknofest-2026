magic
tech sky130A
magscale 1 2
timestamp 1771116256
<< nwell >>
rect -1399 -528 1399 528
<< pmos >>
rect -1203 -308 -953 380
rect -895 -308 -645 380
rect -587 -308 -337 380
rect -279 -308 -29 380
rect 29 -308 279 380
rect 337 -308 587 380
rect 645 -308 895 380
rect 953 -308 1203 380
<< pdiff >>
rect -1261 368 -1203 380
rect -1261 -296 -1249 368
rect -1215 -296 -1203 368
rect -1261 -308 -1203 -296
rect -953 368 -895 380
rect -953 -296 -941 368
rect -907 -296 -895 368
rect -953 -308 -895 -296
rect -645 368 -587 380
rect -645 -296 -633 368
rect -599 -296 -587 368
rect -645 -308 -587 -296
rect -337 368 -279 380
rect -337 -296 -325 368
rect -291 -296 -279 368
rect -337 -308 -279 -296
rect -29 368 29 380
rect -29 -296 -17 368
rect 17 -296 29 368
rect -29 -308 29 -296
rect 279 368 337 380
rect 279 -296 291 368
rect 325 -296 337 368
rect 279 -308 337 -296
rect 587 368 645 380
rect 587 -296 599 368
rect 633 -296 645 368
rect 587 -308 645 -296
rect 895 368 953 380
rect 895 -296 907 368
rect 941 -296 953 368
rect 895 -308 953 -296
rect 1203 368 1261 380
rect 1203 -296 1215 368
rect 1249 -296 1261 368
rect 1203 -308 1261 -296
<< pdiffc >>
rect -1249 -296 -1215 368
rect -941 -296 -907 368
rect -633 -296 -599 368
rect -325 -296 -291 368
rect -17 -296 17 368
rect 291 -296 325 368
rect 599 -296 633 368
rect 907 -296 941 368
rect 1215 -296 1249 368
<< nsubdiff >>
rect -1363 458 -1267 492
rect 1267 458 1363 492
rect -1363 395 -1329 458
rect 1329 395 1363 458
rect -1363 -458 -1329 -395
rect 1329 -458 1363 -395
rect -1363 -492 -1267 -458
rect 1267 -492 1363 -458
<< nsubdiffcont >>
rect -1267 458 1267 492
rect -1363 -395 -1329 395
rect 1329 -395 1363 395
rect -1267 -492 1267 -458
<< poly >>
rect -1203 380 -953 406
rect -895 380 -645 406
rect -587 380 -337 406
rect -279 380 -29 406
rect 29 380 279 406
rect 337 380 587 406
rect 645 380 895 406
rect 953 380 1203 406
rect -1203 -355 -953 -308
rect -1203 -389 -1187 -355
rect -969 -389 -953 -355
rect -1203 -405 -953 -389
rect -895 -355 -645 -308
rect -895 -389 -879 -355
rect -661 -389 -645 -355
rect -895 -405 -645 -389
rect -587 -355 -337 -308
rect -587 -389 -571 -355
rect -353 -389 -337 -355
rect -587 -405 -337 -389
rect -279 -355 -29 -308
rect -279 -389 -263 -355
rect -45 -389 -29 -355
rect -279 -405 -29 -389
rect 29 -355 279 -308
rect 29 -389 45 -355
rect 263 -389 279 -355
rect 29 -405 279 -389
rect 337 -355 587 -308
rect 337 -389 353 -355
rect 571 -389 587 -355
rect 337 -405 587 -389
rect 645 -355 895 -308
rect 645 -389 661 -355
rect 879 -389 895 -355
rect 645 -405 895 -389
rect 953 -355 1203 -308
rect 953 -389 969 -355
rect 1187 -389 1203 -355
rect 953 -405 1203 -389
<< polycont >>
rect -1187 -389 -969 -355
rect -879 -389 -661 -355
rect -571 -389 -353 -355
rect -263 -389 -45 -355
rect 45 -389 263 -355
rect 353 -389 571 -355
rect 661 -389 879 -355
rect 969 -389 1187 -355
<< locali >>
rect -1363 458 -1267 492
rect 1267 458 1363 492
rect -1363 395 -1329 458
rect 1329 395 1363 458
rect -1249 368 -1215 384
rect -1249 -312 -1215 -296
rect -941 368 -907 384
rect -941 -312 -907 -296
rect -633 368 -599 384
rect -633 -312 -599 -296
rect -325 368 -291 384
rect -325 -312 -291 -296
rect -17 368 17 384
rect -17 -312 17 -296
rect 291 368 325 384
rect 291 -312 325 -296
rect 599 368 633 384
rect 599 -312 633 -296
rect 907 368 941 384
rect 907 -312 941 -296
rect 1215 368 1249 384
rect 1215 -312 1249 -296
rect -1203 -389 -1187 -355
rect -969 -389 -953 -355
rect -895 -389 -879 -355
rect -661 -389 -645 -355
rect -587 -389 -571 -355
rect -353 -389 -337 -355
rect -279 -389 -263 -355
rect -45 -389 -29 -355
rect 29 -389 45 -355
rect 263 -389 279 -355
rect 337 -389 353 -355
rect 571 -389 587 -355
rect 645 -389 661 -355
rect 879 -389 895 -355
rect 953 -389 969 -355
rect 1187 -389 1203 -355
rect -1363 -458 -1329 -395
rect 1329 -458 1363 -395
rect -1363 -492 -1267 -458
rect 1267 -492 1363 -458
<< viali >>
rect -1249 -296 -1215 368
rect -941 -296 -907 368
rect -633 -296 -599 368
rect -325 -296 -291 368
rect -17 -296 17 368
rect 291 -296 325 368
rect 599 -296 633 368
rect 907 -296 941 368
rect 1215 -296 1249 368
rect -1187 -389 -969 -355
rect -879 -389 -661 -355
rect -571 -389 -353 -355
rect -263 -389 -45 -355
rect 45 -389 263 -355
rect 353 -389 571 -355
rect 661 -389 879 -355
rect 969 -389 1187 -355
<< metal1 >>
rect -1255 368 -1209 380
rect -1255 -296 -1249 368
rect -1215 -296 -1209 368
rect -1255 -308 -1209 -296
rect -947 368 -901 380
rect -947 -296 -941 368
rect -907 -296 -901 368
rect -947 -308 -901 -296
rect -639 368 -593 380
rect -639 -296 -633 368
rect -599 -296 -593 368
rect -639 -308 -593 -296
rect -331 368 -285 380
rect -331 -296 -325 368
rect -291 -296 -285 368
rect -331 -308 -285 -296
rect -23 368 23 380
rect -23 -296 -17 368
rect 17 -296 23 368
rect -23 -308 23 -296
rect 285 368 331 380
rect 285 -296 291 368
rect 325 -296 331 368
rect 285 -308 331 -296
rect 593 368 639 380
rect 593 -296 599 368
rect 633 -296 639 368
rect 593 -308 639 -296
rect 901 368 947 380
rect 901 -296 907 368
rect 941 -296 947 368
rect 901 -308 947 -296
rect 1209 368 1255 380
rect 1209 -296 1215 368
rect 1249 -296 1255 368
rect 1209 -308 1255 -296
rect -1199 -355 -957 -349
rect -1199 -389 -1187 -355
rect -969 -389 -957 -355
rect -1199 -395 -957 -389
rect -891 -355 -649 -349
rect -891 -389 -879 -355
rect -661 -389 -649 -355
rect -891 -395 -649 -389
rect -583 -355 -341 -349
rect -583 -389 -571 -355
rect -353 -389 -341 -355
rect -583 -395 -341 -389
rect -275 -355 -33 -349
rect -275 -389 -263 -355
rect -45 -389 -33 -355
rect -275 -395 -33 -389
rect 33 -355 275 -349
rect 33 -389 45 -355
rect 263 -389 275 -355
rect 33 -395 275 -389
rect 341 -355 583 -349
rect 341 -389 353 -355
rect 571 -389 583 -355
rect 341 -395 583 -389
rect 649 -355 891 -349
rect 649 -389 661 -355
rect 879 -389 891 -355
rect 649 -395 891 -389
rect 957 -355 1199 -349
rect 957 -389 969 -355
rect 1187 -389 1199 -355
rect 957 -395 1199 -389
<< properties >>
string FIXED_BBOX -1346 -475 1346 475
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 3.4375 l 1.25 m 1 nf 8 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 class mosfet compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1770979109
<< nmos >>
rect -2087 -531 -1087 469
rect -1029 -531 -29 469
rect 29 -531 1029 469
rect 1087 -531 2087 469
<< ndiff >>
rect -2145 457 -2087 469
rect -2145 -519 -2133 457
rect -2099 -519 -2087 457
rect -2145 -531 -2087 -519
rect -1087 457 -1029 469
rect -1087 -519 -1075 457
rect -1041 -519 -1029 457
rect -1087 -531 -1029 -519
rect -29 457 29 469
rect -29 -519 -17 457
rect 17 -519 29 457
rect -29 -531 29 -519
rect 1029 457 1087 469
rect 1029 -519 1041 457
rect 1075 -519 1087 457
rect 1029 -531 1087 -519
rect 2087 457 2145 469
rect 2087 -519 2099 457
rect 2133 -519 2145 457
rect 2087 -531 2145 -519
<< ndiffc >>
rect -2133 -519 -2099 457
rect -1075 -519 -1041 457
rect -17 -519 17 457
rect 1041 -519 1075 457
rect 2099 -519 2133 457
<< poly >>
rect -2087 541 -1087 557
rect -2087 507 -2071 541
rect -1103 507 -1087 541
rect -2087 469 -1087 507
rect -1029 541 -29 557
rect -1029 507 -1013 541
rect -45 507 -29 541
rect -1029 469 -29 507
rect 29 541 1029 557
rect 29 507 45 541
rect 1013 507 1029 541
rect 29 469 1029 507
rect 1087 541 2087 557
rect 1087 507 1103 541
rect 2071 507 2087 541
rect 1087 469 2087 507
rect -2087 -557 -1087 -531
rect -1029 -557 -29 -531
rect 29 -557 1029 -531
rect 1087 -557 2087 -531
<< polycont >>
rect -2071 507 -1103 541
rect -1013 507 -45 541
rect 45 507 1013 541
rect 1103 507 2071 541
<< locali >>
rect -2087 507 -2071 541
rect -1103 507 -1087 541
rect -1029 507 -1013 541
rect -45 507 -29 541
rect 29 507 45 541
rect 1013 507 1029 541
rect 1087 507 1103 541
rect 2071 507 2087 541
rect -2133 457 -2099 473
rect -2133 -535 -2099 -519
rect -1075 457 -1041 473
rect -1075 -535 -1041 -519
rect -17 457 17 473
rect -17 -535 17 -519
rect 1041 457 1075 473
rect 1041 -535 1075 -519
rect 2099 457 2133 473
rect 2099 -535 2133 -519
<< viali >>
rect -2071 507 -1103 541
rect -1013 507 -45 541
rect 45 507 1013 541
rect 1103 507 2071 541
rect -2133 -519 -2099 457
rect -1075 -519 -1041 457
rect -17 -519 17 457
rect 1041 -519 1075 457
rect 2099 -519 2133 457
<< metal1 >>
rect -2083 541 -1091 547
rect -2083 507 -2071 541
rect -1103 507 -1091 541
rect -2083 501 -1091 507
rect -1025 541 -33 547
rect -1025 507 -1013 541
rect -45 507 -33 541
rect -1025 501 -33 507
rect 33 541 1025 547
rect 33 507 45 541
rect 1013 507 1025 541
rect 33 501 1025 507
rect 1091 541 2083 547
rect 1091 507 1103 541
rect 2071 507 2083 541
rect 1091 501 2083 507
rect -2139 457 -2093 469
rect -2139 -519 -2133 457
rect -2099 -519 -2093 457
rect -2139 -531 -2093 -519
rect -1081 457 -1035 469
rect -1081 -519 -1075 457
rect -1041 -519 -1035 457
rect -1081 -531 -1035 -519
rect -23 457 23 469
rect -23 -519 -17 457
rect 17 -519 23 457
rect -23 -531 23 -519
rect 1035 457 1081 469
rect 1035 -519 1041 457
rect 1075 -519 1081 457
rect 1035 -531 1081 -519
rect 2093 457 2139 469
rect 2093 -519 2099 457
rect 2133 -519 2139 457
rect 2093 -531 2139 -519
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 5.0 l 5.0 m 1 nf 4 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 class mosfet compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1770979109
<< nwell >>
rect -2181 -789 2181 823
<< pmos >>
rect -2087 -689 -1087 761
rect -1029 -689 -29 761
rect 29 -689 1029 761
rect 1087 -689 2087 761
<< pdiff >>
rect -2145 749 -2087 761
rect -2145 -677 -2133 749
rect -2099 -677 -2087 749
rect -2145 -689 -2087 -677
rect -1087 749 -1029 761
rect -1087 -677 -1075 749
rect -1041 -677 -1029 749
rect -1087 -689 -1029 -677
rect -29 749 29 761
rect -29 -677 -17 749
rect 17 -677 29 749
rect -29 -689 29 -677
rect 1029 749 1087 761
rect 1029 -677 1041 749
rect 1075 -677 1087 749
rect 1029 -689 1087 -677
rect 2087 749 2145 761
rect 2087 -677 2099 749
rect 2133 -677 2145 749
rect 2087 -689 2145 -677
<< pdiffc >>
rect -2133 -677 -2099 749
rect -1075 -677 -1041 749
rect -17 -677 17 749
rect 1041 -677 1075 749
rect 2099 -677 2133 749
<< poly >>
rect -2087 761 -1087 787
rect -1029 761 -29 787
rect 29 761 1029 787
rect 1087 761 2087 787
rect -2087 -736 -1087 -689
rect -2087 -770 -2071 -736
rect -1103 -770 -1087 -736
rect -2087 -786 -1087 -770
rect -1029 -736 -29 -689
rect -1029 -770 -1013 -736
rect -45 -770 -29 -736
rect -1029 -786 -29 -770
rect 29 -736 1029 -689
rect 29 -770 45 -736
rect 1013 -770 1029 -736
rect 29 -786 1029 -770
rect 1087 -736 2087 -689
rect 1087 -770 1103 -736
rect 2071 -770 2087 -736
rect 1087 -786 2087 -770
<< polycont >>
rect -2071 -770 -1103 -736
rect -1013 -770 -45 -736
rect 45 -770 1013 -736
rect 1103 -770 2071 -736
<< locali >>
rect -2133 749 -2099 765
rect -2133 -693 -2099 -677
rect -1075 749 -1041 765
rect -1075 -693 -1041 -677
rect -17 749 17 765
rect -17 -693 17 -677
rect 1041 749 1075 765
rect 1041 -693 1075 -677
rect 2099 749 2133 765
rect 2099 -693 2133 -677
rect -2087 -770 -2071 -736
rect -1103 -770 -1087 -736
rect -1029 -770 -1013 -736
rect -45 -770 -29 -736
rect 29 -770 45 -736
rect 1013 -770 1029 -736
rect 1087 -770 1103 -736
rect 2071 -770 2087 -736
<< viali >>
rect -2133 -677 -2099 749
rect -1075 -677 -1041 749
rect -17 -677 17 749
rect 1041 -677 1075 749
rect 2099 -677 2133 749
rect -2071 -770 -1103 -736
rect -1013 -770 -45 -736
rect 45 -770 1013 -736
rect 1103 -770 2071 -736
<< metal1 >>
rect -2139 749 -2093 761
rect -2139 -677 -2133 749
rect -2099 -677 -2093 749
rect -2139 -689 -2093 -677
rect -1081 749 -1035 761
rect -1081 -677 -1075 749
rect -1041 -677 -1035 749
rect -1081 -689 -1035 -677
rect -23 749 23 761
rect -23 -677 -17 749
rect 17 -677 23 749
rect -23 -689 23 -677
rect 1035 749 1081 761
rect 1035 -677 1041 749
rect 1075 -677 1081 749
rect 1035 -689 1081 -677
rect 2093 749 2139 761
rect 2093 -677 2099 749
rect 2133 -677 2139 749
rect 2093 -689 2139 -677
rect -2083 -736 -1091 -730
rect -2083 -770 -2071 -736
rect -1103 -770 -1091 -736
rect -2083 -776 -1091 -770
rect -1025 -736 -33 -730
rect -1025 -770 -1013 -736
rect -45 -770 -33 -736
rect -1025 -776 -33 -770
rect 33 -736 1025 -730
rect 33 -770 45 -736
rect 1013 -770 1025 -736
rect 33 -776 1025 -770
rect 1091 -736 2083 -730
rect 1091 -770 1103 -736
rect 2071 -770 2083 -736
rect 1091 -776 2083 -770
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 7.25 l 5.0 m 1 nf 4 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 class mosfet compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

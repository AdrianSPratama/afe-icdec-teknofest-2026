magic
tech sky130A
magscale 1 2
timestamp 1770979109
<< locali >>
rect -100 410 100 467
rect -100 -467 100 -410
<< rlocali >>
rect -100 -410 100 410
<< properties >>
string gencell sky130_fd_pr__res_generic_l1
string library sky130
string parameters w 1.0 l 4.1 m 1 nx 1 wmin 0.17 lmin 0.17 class resistor rho 12.8 val 52.48 dummy 0 dw 0.0 term 0.0 snake 0 roverlap 0
<< end >>

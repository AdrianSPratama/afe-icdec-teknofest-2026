magic
tech sky130A
magscale 1 2
timestamp 1771413069
<< nwell >>
rect -783 -489 783 489
<< pmos >>
rect -587 -270 -337 270
rect -279 -270 -29 270
rect 29 -270 279 270
rect 337 -270 587 270
<< pdiff >>
rect -645 258 -587 270
rect -645 -258 -633 258
rect -599 -258 -587 258
rect -645 -270 -587 -258
rect -337 258 -279 270
rect -337 -258 -325 258
rect -291 -258 -279 258
rect -337 -270 -279 -258
rect -29 258 29 270
rect -29 -258 -17 258
rect 17 -258 29 258
rect -29 -270 29 -258
rect 279 258 337 270
rect 279 -258 291 258
rect 325 -258 337 258
rect 279 -270 337 -258
rect 587 258 645 270
rect 587 -258 599 258
rect 633 -258 645 258
rect 587 -270 645 -258
<< pdiffc >>
rect -633 -258 -599 258
rect -325 -258 -291 258
rect -17 -258 17 258
rect 291 -258 325 258
rect 599 -258 633 258
<< nsubdiff >>
rect -747 419 -651 453
rect 651 419 747 453
rect -747 357 -713 419
rect 713 357 747 419
rect -747 -419 -713 -357
rect 713 -419 747 -357
rect -747 -453 -651 -419
rect 651 -453 747 -419
<< nsubdiffcont >>
rect -651 419 651 453
rect -747 -357 -713 357
rect 713 -357 747 357
rect -651 -453 651 -419
<< poly >>
rect -587 351 -337 367
rect -587 317 -571 351
rect -353 317 -337 351
rect -587 270 -337 317
rect -279 351 -29 367
rect -279 317 -263 351
rect -45 317 -29 351
rect -279 270 -29 317
rect 29 351 279 367
rect 29 317 45 351
rect 263 317 279 351
rect 29 270 279 317
rect 337 351 587 367
rect 337 317 353 351
rect 571 317 587 351
rect 337 270 587 317
rect -587 -317 -337 -270
rect -587 -351 -571 -317
rect -353 -351 -337 -317
rect -587 -367 -337 -351
rect -279 -317 -29 -270
rect -279 -351 -263 -317
rect -45 -351 -29 -317
rect -279 -367 -29 -351
rect 29 -317 279 -270
rect 29 -351 45 -317
rect 263 -351 279 -317
rect 29 -367 279 -351
rect 337 -317 587 -270
rect 337 -351 353 -317
rect 571 -351 587 -317
rect 337 -367 587 -351
<< polycont >>
rect -571 317 -353 351
rect -263 317 -45 351
rect 45 317 263 351
rect 353 317 571 351
rect -571 -351 -353 -317
rect -263 -351 -45 -317
rect 45 -351 263 -317
rect 353 -351 571 -317
<< locali >>
rect -747 419 -651 453
rect 651 419 747 453
rect -747 357 -713 419
rect 713 357 747 419
rect -587 317 -571 351
rect -353 317 -337 351
rect -279 317 -263 351
rect -45 317 -29 351
rect 29 317 45 351
rect 263 317 279 351
rect 337 317 353 351
rect 571 317 587 351
rect -633 258 -599 274
rect -633 -274 -599 -258
rect -325 258 -291 274
rect -325 -274 -291 -258
rect -17 258 17 274
rect -17 -274 17 -258
rect 291 258 325 274
rect 291 -274 325 -258
rect 599 258 633 274
rect 599 -274 633 -258
rect -587 -351 -571 -317
rect -353 -351 -337 -317
rect -279 -351 -263 -317
rect -45 -351 -29 -317
rect 29 -351 45 -317
rect 263 -351 279 -317
rect 337 -351 353 -317
rect 571 -351 587 -317
rect -747 -419 -713 -357
rect 713 -419 747 -357
rect -747 -453 -651 -419
rect 651 -453 747 -419
<< viali >>
rect -571 317 -353 351
rect -263 317 -45 351
rect 45 317 263 351
rect 353 317 571 351
rect -633 -258 -599 258
rect -325 -258 -291 258
rect -17 -258 17 258
rect 291 -258 325 258
rect 599 -258 633 258
rect -571 -351 -353 -317
rect -263 -351 -45 -317
rect 45 -351 263 -317
rect 353 -351 571 -317
<< metal1 >>
rect -583 351 -341 357
rect -583 317 -571 351
rect -353 317 -341 351
rect -583 311 -341 317
rect -275 351 -33 357
rect -275 317 -263 351
rect -45 317 -33 351
rect -275 311 -33 317
rect 33 351 275 357
rect 33 317 45 351
rect 263 317 275 351
rect 33 311 275 317
rect 341 351 583 357
rect 341 317 353 351
rect 571 317 583 351
rect 341 311 583 317
rect -639 258 -593 270
rect -639 -258 -633 258
rect -599 -258 -593 258
rect -639 -270 -593 -258
rect -331 258 -285 270
rect -331 -258 -325 258
rect -291 -258 -285 258
rect -331 -270 -285 -258
rect -23 258 23 270
rect -23 -258 -17 258
rect 17 -258 23 258
rect -23 -270 23 -258
rect 285 258 331 270
rect 285 -258 291 258
rect 325 -258 331 258
rect 285 -270 331 -258
rect 593 258 639 270
rect 593 -258 599 258
rect 633 -258 639 258
rect 593 -270 639 -258
rect -583 -317 -341 -311
rect -583 -351 -571 -317
rect -353 -351 -341 -317
rect -583 -357 -341 -351
rect -275 -317 -33 -311
rect -275 -351 -263 -317
rect -45 -351 -33 -317
rect -275 -357 -33 -351
rect 33 -317 275 -311
rect 33 -351 45 -317
rect 263 -351 275 -317
rect 33 -357 275 -351
rect 341 -317 583 -311
rect 341 -351 353 -317
rect 571 -351 583 -317
rect 341 -357 583 -351
<< properties >>
string FIXED_BBOX -730 -436 730 436
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 2.7 l 1.25 m 1 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 class mosfet compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

* NGSPICE file created from current-mode-bgr_schematics.ext - technology: sky130A

.subckt sky130_fd_pr__nfet_01v8_RX9YJP a_n73_n100# a_n33_n188# a_15_n100# VSUBS
X0 a_15_n100# a_n33_n188# a_n73_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
C0 a_n33_n188# a_n73_n100# 0.02545f
C1 a_15_n100# a_n73_n100# 0.16211f
C2 a_15_n100# a_n33_n188# 0.02545f
C3 a_15_n100# VSUBS 0.11273f
C4 a_n73_n100# VSUBS 0.11273f
C5 a_n33_n188# VSUBS 0.31312f
.ends

.subckt sky130_fd_pr__res_generic_l1_58A49Y li_n100_n410# li_n100_410# li_n100_n467#
+ VSUBS
R0 li_n100_410# li_n100_n467# sky130_fd_pr__res_generic_l1 w=1 l=4.1
C0 li_n100_n467# VSUBS 0.07444f
C1 li_n100_n410# VSUBS 0.4854f
C2 li_n100_410# VSUBS 0.07444f
.ends

.subckt sky130_fd_pr__res_xhigh_po_1p41_CGMGNJ a_n141_n557# a_n141_125# VSUBS
X0 a_n141_125# a_n141_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
C0 a_n141_n557# a_n141_125# 0.06364f
C1 a_n141_n557# VSUBS 0.77135f
C2 a_n141_125# VSUBS 0.77135f
.ends

.subckt sky130_fd_pr__nfet_01v8_CEKAWC a_n1029_n557# a_1029_n531# a_n2087_n557# a_1087_n557#
+ a_2087_n531# a_n29_n531# a_n1087_n531# a_n2145_n531# a_29_n557# VSUBS
X0 a_1029_n531# a_29_n557# a_n29_n531# VSUBS sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=5
X1 a_n29_n531# a_n1029_n557# a_n1087_n531# VSUBS sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=5
X2 a_2087_n531# a_1087_n557# a_1029_n531# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=5
X3 a_n1087_n531# a_n2087_n557# a_n2145_n531# VSUBS sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=5
C0 a_n2145_n531# a_n1087_n531# 0.06632f
C1 a_n2145_n531# a_n2087_n557# 0.20447f
C2 a_n29_n531# a_n1087_n531# 0.06632f
C3 a_n29_n531# a_1029_n531# 0.06632f
C4 a_n29_n531# a_n1029_n557# 0.20447f
C5 a_n1029_n557# a_n1087_n531# 0.20447f
C6 a_n2087_n557# a_n1087_n531# 0.20447f
C7 a_1029_n531# a_1087_n557# 0.20447f
C8 a_n2087_n557# a_n1029_n557# 0.05942f
C9 a_n29_n531# a_29_n557# 0.20447f
C10 a_1029_n531# a_2087_n531# 0.06632f
C11 a_2087_n531# a_1087_n557# 0.20447f
C12 a_1029_n531# a_29_n557# 0.20447f
C13 a_29_n557# a_1087_n557# 0.05942f
C14 a_29_n557# a_n1029_n557# 0.05942f
C15 a_2087_n531# VSUBS 0.59153f
C16 a_1029_n531# VSUBS 0.3387f
C17 a_n29_n531# VSUBS 0.3387f
C18 a_n1087_n531# VSUBS 0.3387f
C19 a_n2145_n531# VSUBS 0.59153f
C20 a_1087_n557# VSUBS 2.11257f
C21 a_29_n557# VSUBS 2.07776f
C22 a_n1029_n557# VSUBS 2.07776f
C23 a_n2087_n557# VSUBS 2.11257f
.ends

.subckt sky130_fd_pr__pfet_01v8_WYTN36 a_3203_n561# a_n3203_n464# w_n4297_n564# a_1029_n464#
+ a_n4261_n464# a_29_n561# a_2087_n464# a_n1029_n561# a_n29_n464# a_3145_n464# a_n2087_n561#
+ a_1087_n561# a_n1087_n464# a_4203_n464# a_n3145_n561# a_2145_n561# a_n2145_n464#
+ a_n4203_n561# VSUBS
X0 a_n1087_n464# a_n2087_n561# a_n2145_n464# w_n4297_n564# sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=5
X1 a_3145_n464# a_2145_n561# a_2087_n464# w_n4297_n564# sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=5
X2 a_1029_n464# a_29_n561# a_n29_n464# w_n4297_n564# sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=5
X3 a_n2145_n464# a_n3145_n561# a_n3203_n464# w_n4297_n564# sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=5
X4 a_n29_n464# a_n1029_n561# a_n1087_n464# w_n4297_n564# sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=5
X5 a_4203_n464# a_3203_n561# a_3145_n464# w_n4297_n564# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=5
X6 a_n3203_n464# a_n4203_n561# a_n4261_n464# w_n4297_n564# sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=5
X7 a_2087_n464# a_1087_n561# a_1029_n464# w_n4297_n564# sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=5
C0 a_2145_n561# a_3203_n561# 0.0619f
C1 a_n3203_n464# a_n2145_n464# 0.06632f
C2 a_1029_n464# a_1087_n561# 0.20447f
C3 a_2087_n464# a_2145_n561# 0.20447f
C4 a_n1029_n561# a_n1087_n464# 0.20447f
C5 a_n4203_n561# a_n3145_n561# 0.0619f
C6 a_n1087_n464# w_n4297_n564# 0.00513f
C7 a_4203_n464# a_3203_n561# 0.20447f
C8 a_n4203_n561# w_n4297_n564# 0.43217f
C9 a_29_n561# a_n29_n464# 0.20447f
C10 a_3203_n561# w_n4297_n564# 0.43217f
C11 a_2145_n561# w_n4297_n564# 0.42607f
C12 a_n2145_n464# a_n1087_n464# 0.06632f
C13 a_29_n561# a_1087_n561# 0.0619f
C14 a_n4261_n464# w_n4297_n564# 0.01761f
C15 a_29_n561# a_1029_n464# 0.20447f
C16 a_n2087_n561# a_n3145_n561# 0.0619f
C17 a_2087_n464# w_n4297_n564# 0.00513f
C18 a_n2087_n561# a_n1029_n561# 0.0619f
C19 a_n2087_n561# w_n4297_n564# 0.42607f
C20 a_4203_n464# w_n4297_n564# 0.01761f
C21 a_n1087_n464# a_n29_n464# 0.06632f
C22 w_n4297_n564# a_n3145_n561# 0.42607f
C23 a_n1029_n561# w_n4297_n564# 0.42607f
C24 a_n2087_n561# a_n2145_n464# 0.20447f
C25 a_n2145_n464# a_n3145_n561# 0.20447f
C26 a_2145_n561# a_1087_n561# 0.0619f
C27 a_n2145_n464# w_n4297_n564# 0.00513f
C28 a_2087_n464# a_1087_n561# 0.20447f
C29 a_1029_n464# a_2087_n464# 0.06632f
C30 a_3145_n464# a_3203_n561# 0.20447f
C31 a_3145_n464# a_2145_n561# 0.20447f
C32 a_n1029_n561# a_n29_n464# 0.20447f
C33 a_n3203_n464# a_n4203_n561# 0.20447f
C34 a_n29_n464# w_n4297_n564# 0.00513f
C35 a_2087_n464# a_3145_n464# 0.06632f
C36 w_n4297_n564# a_1087_n561# 0.42607f
C37 a_1029_n464# w_n4297_n564# 0.00513f
C38 a_3145_n464# a_4203_n464# 0.06632f
C39 a_n4261_n464# a_n3203_n464# 0.06632f
C40 a_3145_n464# w_n4297_n564# 0.00513f
C41 a_n3203_n464# a_n3145_n561# 0.20447f
C42 a_n3203_n464# w_n4297_n564# 0.00513f
C43 a_n1029_n561# a_29_n561# 0.0619f
C44 a_29_n561# w_n4297_n564# 0.42607f
C45 a_n29_n464# a_1029_n464# 0.06632f
C46 a_n4261_n464# a_n4203_n561# 0.20447f
C47 a_n2087_n561# a_n1087_n464# 0.20447f
C48 a_4203_n464# VSUBS 0.57392f
C49 a_3145_n464# VSUBS 0.33357f
C50 a_2087_n464# VSUBS 0.33357f
C51 a_1029_n464# VSUBS 0.33357f
C52 a_n29_n464# VSUBS 0.33357f
C53 a_n1087_n464# VSUBS 0.33357f
C54 a_n2145_n464# VSUBS 0.33357f
C55 a_n3203_n464# VSUBS 0.33357f
C56 a_n4261_n464# VSUBS 0.57392f
C57 a_3203_n561# VSUBS 1.70728f
C58 a_2145_n561# VSUBS 1.67696f
C59 a_1087_n561# VSUBS 1.67696f
C60 a_29_n561# VSUBS 1.67696f
C61 a_n1029_n561# VSUBS 1.67696f
C62 a_n2087_n561# VSUBS 1.67696f
C63 a_n3145_n561# VSUBS 1.67696f
C64 a_n4203_n561# VSUBS 1.70728f
C65 w_n4297_n564# VSUBS 29.9587f
.ends

.subckt sky130_fd_pr__pfet_01v8_Y44983 a_n73_n100# a_15_n100# w_n109_n200# a_n33_n197#
+ VSUBS
X0 a_15_n100# a_n33_n197# a_n73_n100# w_n109_n200# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
C0 w_n109_n200# a_n33_n197# 0.1045f
C1 w_n109_n200# a_n73_n100# 0.00833f
C2 a_n33_n197# a_15_n100# 0.02364f
C3 a_n73_n100# a_15_n100# 0.16211f
C4 a_n33_n197# a_n73_n100# 0.02364f
C5 w_n109_n200# a_15_n100# 0.00833f
C6 a_15_n100# VSUBS 0.1045f
C7 a_n73_n100# VSUBS 0.1045f
C8 a_n33_n197# VSUBS 0.22112f
C9 w_n109_n200# VSUBS 0.2616f
.ends

.subckt sky130_fd_pr__pfet_01v8_AW5DE3 a_687_n536# a_n387_n536# a_29_n562# w_n781_n598#
+ a_329_n536# a_n687_n562# a_n29_n536# a_n745_n536# a_n329_n562# a_387_n562# VSUBS
X0 a_n387_n536# a_n687_n562# a_n745_n536# w_n781_n598# sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=1.5
X1 a_n29_n536# a_n329_n562# a_n387_n536# w_n781_n598# sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1.5
X2 a_329_n536# a_29_n562# a_n29_n536# w_n781_n598# sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1.5
X3 a_687_n536# a_387_n562# a_329_n536# w_n781_n598# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=1.5
C0 w_n781_n598# a_n745_n536# 0.01762f
C1 a_n29_n536# a_n387_n536# 0.19737f
C2 a_n29_n536# a_29_n562# 0.14205f
C3 a_n387_n536# a_n745_n536# 0.19737f
C4 w_n781_n598# a_n687_n562# 0.15322f
C5 a_387_n562# a_329_n536# 0.14205f
C6 w_n781_n598# a_n329_n562# 0.14711f
C7 a_n387_n536# a_n687_n562# 0.14205f
C8 w_n781_n598# a_387_n562# 0.15322f
C9 a_387_n562# a_687_n536# 0.14205f
C10 a_n687_n562# a_n745_n536# 0.14205f
C11 a_n387_n536# a_n329_n562# 0.14205f
C12 a_n329_n562# a_29_n562# 0.0619f
C13 a_n29_n536# a_n329_n562# 0.14205f
C14 a_29_n562# a_387_n562# 0.0619f
C15 w_n781_n598# a_329_n536# 0.00517f
C16 a_329_n536# a_687_n536# 0.19737f
C17 a_29_n562# a_329_n536# 0.14205f
C18 w_n781_n598# a_687_n536# 0.01762f
C19 a_n29_n536# a_329_n536# 0.19737f
C20 a_n387_n536# w_n781_n598# 0.00517f
C21 a_n687_n562# a_n329_n562# 0.0619f
C22 w_n781_n598# a_29_n562# 0.14711f
C23 a_n29_n536# w_n781_n598# 0.00517f
C24 a_687_n536# VSUBS 0.50929f
C25 a_329_n536# VSUBS 0.20431f
C26 a_n29_n536# VSUBS 0.20431f
C27 a_n387_n536# VSUBS 0.20431f
C28 a_n745_n536# VSUBS 0.50929f
C29 a_387_n562# VSUBS 0.52793f
C30 a_29_n562# VSUBS 0.4976f
C31 a_n329_n562# VSUBS 0.4976f
C32 a_n687_n562# VSUBS 0.52793f
C33 w_n781_n598# VSUBS 5.44513f
.ends

.subckt sky130_fd_pr__pfet_01v8_FX5EQP w_n423_n300# a_n387_n200# a_29_n264# a_329_n200#
+ a_n29_n200# a_n329_n264# VSUBS
X0 a_n29_n200# a_n329_n264# a_n387_n200# w_n423_n300# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=1.5
X1 a_329_n200# a_29_n264# a_n29_n200# w_n423_n300# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=1.5
C0 a_29_n264# a_n29_n200# 0.06051f
C1 w_n423_n300# a_n29_n200# 0.00629f
C2 a_n29_n200# a_329_n200# 0.07938f
C3 a_29_n264# a_n329_n264# 0.07007f
C4 a_n329_n264# w_n423_n300# 0.21995f
C5 a_29_n264# w_n423_n300# 0.21995f
C6 a_29_n264# a_329_n200# 0.06051f
C7 w_n423_n300# a_329_n200# 0.01159f
C8 a_n387_n200# a_n29_n200# 0.07938f
C9 a_n329_n264# a_n387_n200# 0.06051f
C10 w_n423_n300# a_n387_n200# 0.01159f
C11 a_n329_n264# a_n29_n200# 0.06051f
C12 a_329_n200# VSUBS 0.2184f
C13 a_n29_n200# VSUBS 0.09456f
C14 a_n387_n200# VSUBS 0.2184f
C15 a_29_n264# VSUBS 0.52044f
C16 a_n329_n264# VSUBS 0.52044f
C17 w_n423_n300# VSUBS 1.5228f
.ends

.subckt sky130_fd_pr__pfet_01v8_VCUNPM a_500_n349# w_n594_n411# a_n558_n349# a_n500_n375#
+ VSUBS
X0 a_500_n349# a_n500_n375# a_n558_n349# w_n594_n411# sky130_fd_pr__pfet_01v8 ad=0.9077 pd=6.84 as=0.9077 ps=6.84 w=3.13 l=5
C0 a_n558_n349# a_n500_n375# 0.13074f
C1 a_n500_n375# w_n594_n411# 0.43969f
C2 a_n558_n349# w_n594_n411# 0.01314f
C3 a_n500_n375# a_500_n349# 0.13074f
C4 a_n558_n349# a_500_n349# 0.0416f
C5 w_n594_n411# a_500_n349# 0.01314f
C6 a_500_n349# VSUBS 0.36854f
C7 a_n558_n349# VSUBS 0.36854f
C8 a_n500_n375# VSUBS 1.7574f
C9 w_n594_n411# VSUBS 2.80843f
.ends

.subckt sky130_fd_pr__pfet_01v8_MW3DW6 a_n1029_n787# a_1029_n761# a_n29_n761# a_n1087_n761#
+ w_n1123_n823# a_29_n787# VSUBS
X0 a_1029_n761# a_29_n787# a_n29_n761# w_n1123_n823# sky130_fd_pr__pfet_01v8 ad=2.1025 pd=15.08 as=1.05125 ps=7.54 w=7.25 l=5
X1 a_n29_n761# a_n1029_n787# a_n1087_n761# w_n1123_n823# sky130_fd_pr__pfet_01v8 ad=1.05125 pd=7.54 as=2.1025 ps=15.08 w=7.25 l=5
C0 a_29_n787# a_n29_n761# 0.29318f
C1 w_n1123_n823# a_n29_n761# 0.00513f
C2 a_n29_n761# a_1029_n761# 0.09607f
C3 a_29_n787# a_n1029_n787# 0.0619f
C4 a_n1029_n787# w_n1123_n823# 0.43152f
C5 a_29_n787# w_n1123_n823# 0.43152f
C6 a_29_n787# a_1029_n761# 0.29318f
C7 w_n1123_n823# a_1029_n761# 0.02297f
C8 a_n1087_n761# a_n29_n761# 0.09607f
C9 a_n1029_n787# a_n1087_n761# 0.29318f
C10 w_n1123_n823# a_n1087_n761# 0.02297f
C11 a_n1029_n787# a_n29_n761# 0.29318f
C12 a_1029_n761# VSUBS 0.82104f
C13 a_n29_n761# VSUBS 0.47463f
C14 a_n1087_n761# VSUBS 0.82104f
C15 a_29_n787# VSUBS 1.69504f
C16 a_n1029_n787# VSUBS 1.69504f
C17 w_n1123_n823# VSUBS 10.8617f
.ends

.subckt current-mode-bgr_schematics VDD IREF VSS
XXM13 VSS VSS m1_n1020_n1240# VSS sky130_fd_pr__nfet_01v8_RX9YJP
XR1 R9/li_n100_n410# li_3100_120# VSS VSS sky130_fd_pr__res_generic_l1_58A49Y
Xsky130_fd_pr__nfet_01v8_RX9YJP_0 VSS m1_5520_n1460# VSS VSS sky130_fd_pr__nfet_01v8_RX9YJP
XR3 R9/li_n100_n410# li_3100_120# VSS VSS sky130_fd_pr__res_generic_l1_58A49Y
XR4 R9/li_n100_n410# li_3100_120# VSS VSS sky130_fd_pr__res_generic_l1_58A49Y
XR5 R9/li_n100_n410# li_3100_120# VSS VSS sky130_fd_pr__res_generic_l1_58A49Y
XR6 R9/li_n100_n410# li_3100_120# VSS VSS sky130_fd_pr__res_generic_l1_58A49Y
XXR2 m1_2460_n2160# m1_2800_n1480# VSS sky130_fd_pr__res_xhigh_po_1p41_CGMGNJ
XR7 R9/li_n100_n410# li_3100_120# VSS VSS sky130_fd_pr__res_generic_l1_58A49Y
XXR12 m1_3140_n2140# m1_2800_n1480# VSS sky130_fd_pr__res_xhigh_po_1p41_CGMGNJ
XR9 R9/li_n100_n410# li_3100_120# VSS VSS sky130_fd_pr__res_generic_l1_58A49Y
XR8 R9/li_n100_n410# li_3100_120# VSS VSS sky130_fd_pr__res_generic_l1_58A49Y
XXR13 m1_3140_n2140# m1_3480_n1460# VSS sky130_fd_pr__res_xhigh_po_1p41_CGMGNJ
XXR14 m1_3820_n2160# m1_3480_n1460# VSS sky130_fd_pr__res_xhigh_po_1p41_CGMGNJ
XXM1 m1_n200_2800# li_3100_120# m1_n200_2800# m1_n200_2800# m1_n200_2800# m1_n720_1500#
+ VSS m1_n200_2800# m1_n200_2800# VSS sky130_fd_pr__nfet_01v8_CEKAWC
XR10 R9/li_n100_n410# li_3100_120# VSS VSS sky130_fd_pr__res_generic_l1_58A49Y
XXR15 m1_3820_n2160# m1_4160_n1460# VSS sky130_fd_pr__res_xhigh_po_1p41_CGMGNJ
XR21 R9/li_n100_n410# li_3100_120# VSS VSS sky130_fd_pr__res_generic_l1_58A49Y
XXM3 m1_n720_1500# VDD VDD VDD m1_n200_2800# m1_n720_1500# m1_n720_1500# m1_n720_1500#
+ m1_n200_2800# VDD m1_n720_1500# m1_n720_1500# VDD m1_n200_2800# m1_n720_1500# m1_n720_1500#
+ m1_n720_1500# m1_n720_1500# VSS sky130_fd_pr__pfet_01v8_WYTN36
XXR16 m1_4500_n2160# m1_4160_n1460# VSS sky130_fd_pr__res_xhigh_po_1p41_CGMGNJ
XXR17 m1_4500_n2160# m1_4840_n1460# VSS sky130_fd_pr__res_xhigh_po_1p41_CGMGNJ
XXR18 m1_5180_n2140# m1_4840_n1460# VSS sky130_fd_pr__res_xhigh_po_1p41_CGMGNJ
XXM5 VDD m1_n200_2800# VDD VSS VSS sky130_fd_pr__pfet_01v8_Y44983
XXR19 m1_5180_n2140# m1_5520_n1460# VSS sky130_fd_pr__res_xhigh_po_1p41_CGMGNJ
XXM6 m1_640_300# VDD m1_n720_1500# VDD VDD m1_n720_1500# VSS m1_n800_300# m1_n720_1500#
+ m1_n720_1500# VSS sky130_fd_pr__pfet_01v8_AW5DE3
XXM8 VDD m1_n1020_n1240# m1_n1020_n1240# m1_5520_n1460# VDD m1_n1020_n1240# VSS sky130_fd_pr__pfet_01v8_FX5EQP
Xsky130_fd_pr__pfet_01v8_AW5DE3_0 VSS VDD m1_n720_1500# VDD VDD m1_n720_1500# VSS
+ VSS m1_n720_1500# m1_n720_1500# VSS sky130_fd_pr__pfet_01v8_AW5DE3
Xsky130_fd_pr__pfet_01v8_VCUNPM_0 VDD VDD IREF m1_n720_1500# VSS sky130_fd_pr__pfet_01v8_VCUNPM
Xsky130_fd_pr__res_xhigh_po_1p41_CGMGNJ_0 m1_2460_n2160# VSS VSS sky130_fd_pr__res_xhigh_po_1p41_CGMGNJ
Xsky130_fd_pr__pfet_01v8_MW3DW6_0 m1_n1020_n1240# IREF VDD IREF VDD m1_n1020_n1240#
+ VSS sky130_fd_pr__pfet_01v8_MW3DW6
XXM10 IREF VDD VDD m1_n720_1500# VSS sky130_fd_pr__pfet_01v8_VCUNPM
XXM11 m1_n1020_n1240# IREF VDD IREF VDD m1_n1020_n1240# VSS sky130_fd_pr__pfet_01v8_MW3DW6
C0 R9/li_n100_n410# m1_4160_n1460# 0.02448f
C1 m1_4160_n1460# m1_5520_n1460# 0.00125f
C2 m1_640_300# m1_n720_1500# 0.0825f
C3 m1_3480_n1460# m1_n720_1500# 0.00454f
C4 li_3100_120# VDD 0.01501f
C5 m1_4840_n1460# m1_n1020_n1240# 0.25438f
C6 R9/li_n100_n410# m1_n720_1500# 0.0037f
C7 li_3100_120# m1_4160_n1460# 0.00811f
C8 m1_5520_n1460# m1_n720_1500# 0.03916f
C9 m1_3820_n2160# m1_n1020_n1240# 0.03062f
C10 li_3100_120# m1_n720_1500# 1.84338f
C11 m1_2800_n1480# VDD 0
C12 m1_2800_n1480# m1_3140_n2140# 0.00493f
C13 m1_n200_2800# VDD 3.71212f
C14 m1_5180_n2140# m1_n1020_n1240# 0.03049f
C15 m1_5520_n1460# IREF 0.514f
C16 m1_2800_n1480# m1_4160_n1460# 0
C17 m1_4500_n2160# m1_4840_n1460# 0.00259f
C18 m1_4160_n1460# m1_n200_2800# 0
C19 VDD m1_n1020_n1240# 12.79605f
C20 m1_3140_n2140# m1_n1020_n1240# 0.03049f
C21 m1_2800_n1480# m1_2460_n2160# 0.00464f
C22 m1_2800_n1480# m1_n720_1500# 0.00166f
C23 m1_4160_n1460# m1_n1020_n1240# 0.25438f
C24 m1_n800_300# m1_n1020_n1240# 0
C25 m1_n200_2800# m1_n720_1500# 5.6971f
C26 m1_3820_n2160# m1_4500_n2160# 0.43168f
C27 m1_2460_n2160# m1_n1020_n1240# 0.03234f
C28 m1_4500_n2160# m1_5180_n2140# 0.42687f
C29 m1_n720_1500# m1_n1020_n1240# 0.83816f
C30 R9/li_n100_n410# m1_3480_n1460# 0.02448f
C31 m1_n200_2800# IREF 0
C32 m1_4500_n2160# VDD 0.01339f
C33 R9/li_n100_n410# m1_5520_n1460# 0.01279f
C34 m1_3140_n2140# m1_4500_n2160# 0
C35 m1_4160_n1460# m1_4500_n2160# 0.00258f
C36 li_3100_120# m1_3480_n1460# 0.00788f
C37 m1_n1020_n1240# IREF 1.68036f
C38 li_3100_120# R9/li_n100_n410# 0.09702f
C39 m1_4500_n2160# m1_n720_1500# 0.02999f
C40 m1_2800_n1480# m1_3480_n1460# 0.42657f
C41 m1_n200_2800# m1_640_300# 0.05965f
C42 m1_3480_n1460# m1_n200_2800# 0
C43 R9/li_n100_n410# m1_2800_n1480# 0.01238f
C44 R9/li_n100_n410# m1_n200_2800# 0.03076f
C45 m1_4840_n1460# m1_5180_n2140# 0.00287f
C46 m1_640_300# m1_n1020_n1240# 0
C47 m1_n200_2800# m1_5520_n1460# 0.01838f
C48 m1_3480_n1460# m1_n1020_n1240# 0.25459f
C49 m1_4840_n1460# VDD 0
C50 R9/li_n100_n410# m1_n1020_n1240# 0.74858f
C51 li_3100_120# m1_2800_n1480# 0
C52 m1_5520_n1460# m1_n1020_n1240# 3.64118f
C53 li_3100_120# m1_n200_2800# 3.64665f
C54 m1_4160_n1460# m1_4840_n1460# 0.42654f
C55 m1_3820_n2160# m1_5180_n2140# 0
C56 li_3100_120# m1_n1020_n1240# 0.09869f
C57 m1_3820_n2160# VDD 0.01339f
C58 m1_3140_n2140# m1_3820_n2160# 0.42683f
C59 m1_4840_n1460# m1_n720_1500# 0.00164f
C60 m1_3820_n2160# m1_4160_n1460# 0.00259f
C61 m1_5180_n2140# VDD 0.01531f
C62 m1_2800_n1480# m1_n200_2800# 0
C63 m1_3140_n2140# m1_5180_n2140# 0
C64 R9/li_n100_n410# m1_4500_n2160# 0
C65 m1_3820_n2160# m1_2460_n2160# 0
C66 m1_3140_n2140# VDD 0.01264f
C67 m1_3820_n2160# m1_n720_1500# 0.02999f
C68 m1_2800_n1480# m1_n1020_n1240# 0.25703f
C69 m1_4840_n1460# IREF 0
C70 m1_n200_2800# m1_n1020_n1240# 0.08386f
C71 m1_4160_n1460# VDD 0
C72 m1_n800_300# VDD 0.48583f
C73 m1_5180_n2140# m1_n720_1500# 0.02953f
C74 m1_2460_n2160# VDD 0.01673f
C75 m1_3140_n2140# m1_2460_n2160# 0.42687f
C76 m1_n720_1500# VDD 41.32107f
C77 m1_3140_n2140# m1_n720_1500# 0.02953f
C78 m1_4160_n1460# m1_n720_1500# 0.0028f
C79 m1_5180_n2140# IREF 0.01699f
C80 m1_n800_300# m1_n720_1500# 0.10129f
C81 m1_2460_n2160# m1_n720_1500# 0.02999f
C82 VDD IREF 14.17803f
C83 R9/li_n100_n410# m1_4840_n1460# 0.01027f
C84 m1_4500_n2160# m1_n1020_n1240# 0.03062f
C85 m1_4840_n1460# m1_5520_n1460# 0.43295f
C86 m1_3480_n1460# m1_3820_n2160# 0.00258f
C87 m1_2460_n2160# IREF 0.01586f
C88 li_3100_120# m1_4840_n1460# 0.00647f
C89 m1_n720_1500# IREF 2.49635f
C90 R9/li_n100_n410# m1_3820_n2160# 0
C91 m1_640_300# VDD 0.41153f
C92 m1_3480_n1460# VDD 0
C93 m1_5520_n1460# m1_5180_n2140# 0.00287f
C94 m1_3140_n2140# m1_3480_n1460# 0.00287f
C95 m1_3480_n1460# m1_4160_n1460# 0.42654f
C96 m1_2800_n1480# m1_4840_n1460# 0
C97 m1_5520_n1460# VDD 3.91857f
C98 R9/li_n100_n410# m1_3140_n2140# 0
C99 m1_4840_n1460# m1_n200_2800# 0
C100 IREF VSS 3.01077f
C101 m1_n1020_n1240# VSS 9.50681f
C102 VDD VSS 0.21929p
C103 m1_n720_1500# VSS 14.94089f
C104 m1_2460_n2160# VSS 0.73141f
C105 m1_640_300# VSS 0.21166f
C106 m1_n800_300# VSS 0.26131f
C107 m1_5180_n2140# VSS 0.71312f
C108 m1_5520_n1460# VSS 3.73797f
C109 m1_n200_2800# VSS 15.02407f
C110 m1_4840_n1460# VSS 0.57986f
C111 m1_4500_n2160# VSS 0.56819f
C112 m1_4160_n1460# VSS 0.55907f
C113 m1_3820_n2160# VSS 0.56743f
C114 m1_3480_n1460# VSS 0.55797f
C115 m1_3140_n2140# VSS 0.55109f
C116 m1_2800_n1480# VSS 1.01531f
C117 li_3100_120# VSS 2.10081f
C118 R9/li_n100_n410# VSS 2.49061f
.ends


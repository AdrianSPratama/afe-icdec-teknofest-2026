magic
tech sky130A
magscale 1 2
timestamp 1770979109
<< pwell >>
rect -2283 -710 2283 710
<< nmos >>
rect -2087 -500 -1087 500
rect -1029 -500 -29 500
rect 29 -500 1029 500
rect 1087 -500 2087 500
<< ndiff >>
rect -2145 488 -2087 500
rect -2145 -488 -2133 488
rect -2099 -488 -2087 488
rect -2145 -500 -2087 -488
rect -1087 488 -1029 500
rect -1087 -488 -1075 488
rect -1041 -488 -1029 488
rect -1087 -500 -1029 -488
rect -29 488 29 500
rect -29 -488 -17 488
rect 17 -488 29 488
rect -29 -500 29 -488
rect 1029 488 1087 500
rect 1029 -488 1041 488
rect 1075 -488 1087 488
rect 1029 -500 1087 -488
rect 2087 488 2145 500
rect 2087 -488 2099 488
rect 2133 -488 2145 488
rect 2087 -500 2145 -488
<< ndiffc >>
rect -2133 -488 -2099 488
rect -1075 -488 -1041 488
rect -17 -488 17 488
rect 1041 -488 1075 488
rect 2099 -488 2133 488
<< psubdiff >>
rect -2247 640 -2151 674
rect 2151 640 2247 674
rect -2247 578 -2213 640
rect 2213 578 2247 640
rect -2247 -640 -2213 -578
rect 2213 -640 2247 -578
rect -2247 -674 -2151 -640
rect 2151 -674 2247 -640
<< psubdiffcont >>
rect -2151 640 2151 674
rect -2247 -578 -2213 578
rect 2213 -578 2247 578
rect -2151 -674 2151 -640
<< poly >>
rect -2087 572 -1087 588
rect -2087 538 -2071 572
rect -1103 538 -1087 572
rect -2087 500 -1087 538
rect -1029 572 -29 588
rect -1029 538 -1013 572
rect -45 538 -29 572
rect -1029 500 -29 538
rect 29 572 1029 588
rect 29 538 45 572
rect 1013 538 1029 572
rect 29 500 1029 538
rect 1087 572 2087 588
rect 1087 538 1103 572
rect 2071 538 2087 572
rect 1087 500 2087 538
rect -2087 -538 -1087 -500
rect -2087 -572 -2071 -538
rect -1103 -572 -1087 -538
rect -2087 -588 -1087 -572
rect -1029 -538 -29 -500
rect -1029 -572 -1013 -538
rect -45 -572 -29 -538
rect -1029 -588 -29 -572
rect 29 -538 1029 -500
rect 29 -572 45 -538
rect 1013 -572 1029 -538
rect 29 -588 1029 -572
rect 1087 -538 2087 -500
rect 1087 -572 1103 -538
rect 2071 -572 2087 -538
rect 1087 -588 2087 -572
<< polycont >>
rect -2071 538 -1103 572
rect -1013 538 -45 572
rect 45 538 1013 572
rect 1103 538 2071 572
rect -2071 -572 -1103 -538
rect -1013 -572 -45 -538
rect 45 -572 1013 -538
rect 1103 -572 2071 -538
<< locali >>
rect -2247 640 -2151 674
rect 2151 640 2247 674
rect -2247 578 -2213 640
rect 2213 578 2247 640
rect -2087 538 -2071 572
rect -1103 538 -1087 572
rect -1029 538 -1013 572
rect -45 538 -29 572
rect 29 538 45 572
rect 1013 538 1029 572
rect 1087 538 1103 572
rect 2071 538 2087 572
rect -2133 488 -2099 504
rect -2133 -504 -2099 -488
rect -1075 488 -1041 504
rect -1075 -504 -1041 -488
rect -17 488 17 504
rect -17 -504 17 -488
rect 1041 488 1075 504
rect 1041 -504 1075 -488
rect 2099 488 2133 504
rect 2099 -504 2133 -488
rect -2087 -572 -2071 -538
rect -1103 -572 -1087 -538
rect -1029 -572 -1013 -538
rect -45 -572 -29 -538
rect 29 -572 45 -538
rect 1013 -572 1029 -538
rect 1087 -572 1103 -538
rect 2071 -572 2087 -538
rect -2247 -640 -2213 -578
rect 2213 -640 2247 -578
rect -2247 -674 -2151 -640
rect 2151 -674 2247 -640
<< viali >>
rect -2071 538 -1103 572
rect -1013 538 -45 572
rect 45 538 1013 572
rect 1103 538 2071 572
rect -2133 -488 -2099 488
rect -1075 -488 -1041 488
rect -17 -488 17 488
rect 1041 -488 1075 488
rect 2099 -488 2133 488
rect -2071 -572 -1103 -538
rect -1013 -572 -45 -538
rect 45 -572 1013 -538
rect 1103 -572 2071 -538
<< metal1 >>
rect -2083 572 -1091 578
rect -2083 538 -2071 572
rect -1103 538 -1091 572
rect -2083 532 -1091 538
rect -1025 572 -33 578
rect -1025 538 -1013 572
rect -45 538 -33 572
rect -1025 532 -33 538
rect 33 572 1025 578
rect 33 538 45 572
rect 1013 538 1025 572
rect 33 532 1025 538
rect 1091 572 2083 578
rect 1091 538 1103 572
rect 2071 538 2083 572
rect 1091 532 2083 538
rect -2139 488 -2093 500
rect -2139 -488 -2133 488
rect -2099 -488 -2093 488
rect -2139 -500 -2093 -488
rect -1081 488 -1035 500
rect -1081 -488 -1075 488
rect -1041 -488 -1035 488
rect -1081 -500 -1035 -488
rect -23 488 23 500
rect -23 -488 -17 488
rect 17 -488 23 488
rect -23 -500 23 -488
rect 1035 488 1081 500
rect 1035 -488 1041 488
rect 1075 -488 1081 488
rect 1035 -500 1081 -488
rect 2093 488 2139 500
rect 2093 -488 2099 488
rect 2133 -488 2139 488
rect 2093 -500 2139 -488
rect -2083 -538 -1091 -532
rect -2083 -572 -2071 -538
rect -1103 -572 -1091 -538
rect -2083 -578 -1091 -572
rect -1025 -538 -33 -532
rect -1025 -572 -1013 -538
rect -45 -572 -33 -538
rect -1025 -578 -33 -572
rect 33 -538 1025 -532
rect 33 -572 45 -538
rect 1013 -572 1025 -538
rect 33 -578 1025 -572
rect 1091 -538 2083 -532
rect 1091 -572 1103 -538
rect 2071 -572 2083 -538
rect 1091 -578 2083 -572
<< properties >>
string FIXED_BBOX -2230 -657 2230 657
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 5.0 l 5.0 m 1 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 class mosfet compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

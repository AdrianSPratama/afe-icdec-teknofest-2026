magic
tech sky130A
magscale 1 2
timestamp 1771413069
<< pwell >>
rect -783 -479 783 479
<< nmos >>
rect -587 -269 -337 331
rect -279 -269 -29 331
rect 29 -269 279 331
rect 337 -269 587 331
<< ndiff >>
rect -645 319 -587 331
rect -645 -257 -633 319
rect -599 -257 -587 319
rect -645 -269 -587 -257
rect -337 319 -279 331
rect -337 -257 -325 319
rect -291 -257 -279 319
rect -337 -269 -279 -257
rect -29 319 29 331
rect -29 -257 -17 319
rect 17 -257 29 319
rect -29 -269 29 -257
rect 279 319 337 331
rect 279 -257 291 319
rect 325 -257 337 319
rect 279 -269 337 -257
rect 587 319 645 331
rect 587 -257 599 319
rect 633 -257 645 319
rect 587 -269 645 -257
<< ndiffc >>
rect -633 -257 -599 319
rect -325 -257 -291 319
rect -17 -257 17 319
rect 291 -257 325 319
rect 599 -257 633 319
<< psubdiff >>
rect -747 409 -651 443
rect 651 409 747 443
rect -747 347 -713 409
rect 713 347 747 409
rect -747 -409 -713 -347
rect 713 -409 747 -347
rect -747 -443 -651 -409
rect 651 -443 747 -409
<< psubdiffcont >>
rect -651 409 651 443
rect -747 -347 -713 347
rect 713 -347 747 347
rect -651 -443 651 -409
<< poly >>
rect -587 331 -337 357
rect -279 331 -29 357
rect 29 331 279 357
rect 337 331 587 357
rect -587 -307 -337 -269
rect -587 -341 -571 -307
rect -353 -341 -337 -307
rect -587 -357 -337 -341
rect -279 -307 -29 -269
rect -279 -341 -263 -307
rect -45 -341 -29 -307
rect -279 -357 -29 -341
rect 29 -307 279 -269
rect 29 -341 45 -307
rect 263 -341 279 -307
rect 29 -357 279 -341
rect 337 -307 587 -269
rect 337 -341 353 -307
rect 571 -341 587 -307
rect 337 -357 587 -341
<< polycont >>
rect -571 -341 -353 -307
rect -263 -341 -45 -307
rect 45 -341 263 -307
rect 353 -341 571 -307
<< locali >>
rect -747 409 -651 443
rect 651 409 747 443
rect -747 347 -713 409
rect 713 347 747 409
rect -633 319 -599 335
rect -633 -273 -599 -257
rect -325 319 -291 335
rect -325 -273 -291 -257
rect -17 319 17 335
rect -17 -273 17 -257
rect 291 319 325 335
rect 291 -273 325 -257
rect 599 319 633 335
rect 599 -273 633 -257
rect -587 -341 -571 -307
rect -353 -341 -337 -307
rect -279 -341 -263 -307
rect -45 -341 -29 -307
rect 29 -341 45 -307
rect 263 -341 279 -307
rect 337 -341 353 -307
rect 571 -341 587 -307
rect -747 -409 -713 -347
rect 713 -409 747 -347
rect -747 -443 -651 -409
rect 651 -443 747 -409
<< viali >>
rect -633 -257 -599 319
rect -325 -257 -291 319
rect -17 -257 17 319
rect 291 -257 325 319
rect 599 -257 633 319
rect -571 -341 -353 -307
rect -263 -341 -45 -307
rect 45 -341 263 -307
rect 353 -341 571 -307
<< metal1 >>
rect -639 319 -593 331
rect -639 -257 -633 319
rect -599 -257 -593 319
rect -639 -269 -593 -257
rect -331 319 -285 331
rect -331 -257 -325 319
rect -291 -257 -285 319
rect -331 -269 -285 -257
rect -23 319 23 331
rect -23 -257 -17 319
rect 17 -257 23 319
rect -23 -269 23 -257
rect 285 319 331 331
rect 285 -257 291 319
rect 325 -257 331 319
rect 285 -269 331 -257
rect 593 319 639 331
rect 593 -257 599 319
rect 633 -257 639 319
rect 593 -269 639 -257
rect -583 -307 -341 -301
rect -583 -341 -571 -307
rect -353 -341 -341 -307
rect -583 -347 -341 -341
rect -275 -307 -33 -301
rect -275 -341 -263 -307
rect -45 -341 -33 -307
rect -275 -347 -33 -341
rect 33 -307 275 -301
rect 33 -341 45 -307
rect 263 -341 275 -307
rect 33 -347 275 -341
rect 341 -307 583 -301
rect 341 -341 353 -307
rect 571 -341 583 -307
rect 341 -347 583 -341
<< properties >>
string FIXED_BBOX -730 -426 730 426
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 3.0 l 1.25 m 1 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 class mosfet compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

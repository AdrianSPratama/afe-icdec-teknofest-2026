magic
tech sky130A
magscale 1 2
timestamp 1771418038
<< error_p >>
rect -681 1915 681 2166
rect -681 650 681 901
rect -681 -615 681 -364
rect -681 -1880 681 -1629
<< nwell >>
rect -681 1915 681 3177
rect -681 650 681 1912
rect -681 -615 681 647
rect -681 -1880 681 -618
rect -681 -3145 681 -1883
<< pmos >>
rect -587 2015 -337 3115
rect -279 2015 -29 3115
rect 29 2015 279 3115
rect 337 2015 587 3115
rect -587 750 -337 1850
rect -279 750 -29 1850
rect 29 750 279 1850
rect 337 750 587 1850
rect -587 -515 -337 585
rect -279 -515 -29 585
rect 29 -515 279 585
rect 337 -515 587 585
rect -587 -1780 -337 -680
rect -279 -1780 -29 -680
rect 29 -1780 279 -680
rect 337 -1780 587 -680
rect -587 -3045 -337 -1945
rect -279 -3045 -29 -1945
rect 29 -3045 279 -1945
rect 337 -3045 587 -1945
<< pdiff >>
rect -645 2834 -587 3115
rect -645 2296 -633 2834
rect -599 2296 -587 2834
rect -645 2015 -587 2296
rect -337 2834 -279 3115
rect -337 2296 -325 2834
rect -291 2296 -279 2834
rect -337 2015 -279 2296
rect -29 2834 29 3115
rect -29 2296 -17 2834
rect 17 2296 29 2834
rect -29 2015 29 2296
rect 279 2834 337 3115
rect 279 2296 291 2834
rect 325 2296 337 2834
rect 279 2015 337 2296
rect 587 2834 645 3115
rect 587 2296 599 2834
rect 633 2296 645 2834
rect 587 2015 645 2296
rect -645 1569 -587 1850
rect -645 1031 -633 1569
rect -599 1031 -587 1569
rect -645 750 -587 1031
rect -337 1569 -279 1850
rect -337 1031 -325 1569
rect -291 1031 -279 1569
rect -337 750 -279 1031
rect -29 1569 29 1850
rect -29 1031 -17 1569
rect 17 1031 29 1569
rect -29 750 29 1031
rect 279 1569 337 1850
rect 279 1031 291 1569
rect 325 1031 337 1569
rect 279 750 337 1031
rect 587 1569 645 1850
rect 587 1031 599 1569
rect 633 1031 645 1569
rect 587 750 645 1031
rect -645 304 -587 585
rect -645 -234 -633 304
rect -599 -234 -587 304
rect -645 -515 -587 -234
rect -337 304 -279 585
rect -337 -234 -325 304
rect -291 -234 -279 304
rect -337 -515 -279 -234
rect -29 304 29 585
rect -29 -234 -17 304
rect 17 -234 29 304
rect -29 -515 29 -234
rect 279 304 337 585
rect 279 -234 291 304
rect 325 -234 337 304
rect 279 -515 337 -234
rect 587 304 645 585
rect 587 -234 599 304
rect 633 -234 645 304
rect 587 -515 645 -234
rect -645 -961 -587 -680
rect -645 -1499 -633 -961
rect -599 -1499 -587 -961
rect -645 -1780 -587 -1499
rect -337 -961 -279 -680
rect -337 -1499 -325 -961
rect -291 -1499 -279 -961
rect -337 -1780 -279 -1499
rect -29 -961 29 -680
rect -29 -1499 -17 -961
rect 17 -1499 29 -961
rect -29 -1780 29 -1499
rect 279 -961 337 -680
rect 279 -1499 291 -961
rect 325 -1499 337 -961
rect 279 -1780 337 -1499
rect 587 -961 645 -680
rect 587 -1499 599 -961
rect 633 -1499 645 -961
rect 587 -1780 645 -1499
rect -645 -2226 -587 -1945
rect -645 -2764 -633 -2226
rect -599 -2764 -587 -2226
rect -645 -3045 -587 -2764
rect -337 -2226 -279 -1945
rect -337 -2764 -325 -2226
rect -291 -2764 -279 -2226
rect -337 -3045 -279 -2764
rect -29 -2226 29 -1945
rect -29 -2764 -17 -2226
rect 17 -2764 29 -2226
rect -29 -3045 29 -2764
rect 279 -2226 337 -1945
rect 279 -2764 291 -2226
rect 325 -2764 337 -2226
rect 279 -3045 337 -2764
rect 587 -2226 645 -1945
rect 587 -2764 599 -2226
rect 633 -2764 645 -2226
rect 587 -3045 645 -2764
<< pdiffc >>
rect -633 2296 -599 2834
rect -325 2296 -291 2834
rect -17 2296 17 2834
rect 291 2296 325 2834
rect 599 2296 633 2834
rect -633 1031 -599 1569
rect -325 1031 -291 1569
rect -17 1031 17 1569
rect 291 1031 325 1569
rect 599 1031 633 1569
rect -633 -234 -599 304
rect -325 -234 -291 304
rect -17 -234 17 304
rect 291 -234 325 304
rect 599 -234 633 304
rect -633 -1499 -599 -961
rect -325 -1499 -291 -961
rect -17 -1499 17 -961
rect 291 -1499 325 -961
rect 599 -1499 633 -961
rect -633 -2764 -599 -2226
rect -325 -2764 -291 -2226
rect -17 -2764 17 -2226
rect 291 -2764 325 -2226
rect 599 -2764 633 -2226
<< poly >>
rect -587 3115 -337 3141
rect -279 3115 -29 3141
rect 29 3115 279 3141
rect 337 3115 587 3141
rect -587 1968 -337 2015
rect -587 1934 -571 1968
rect -353 1934 -337 1968
rect -587 1918 -337 1934
rect -279 1968 -29 2015
rect -279 1934 -263 1968
rect -45 1934 -29 1968
rect -279 1918 -29 1934
rect 29 1968 279 2015
rect 29 1934 45 1968
rect 263 1934 279 1968
rect 29 1918 279 1934
rect 337 1968 587 2015
rect 337 1934 353 1968
rect 571 1934 587 1968
rect 337 1918 587 1934
rect -587 1850 -337 1876
rect -279 1850 -29 1876
rect 29 1850 279 1876
rect 337 1850 587 1876
rect -587 703 -337 750
rect -587 669 -571 703
rect -353 669 -337 703
rect -587 653 -337 669
rect -279 703 -29 750
rect -279 669 -263 703
rect -45 669 -29 703
rect -279 653 -29 669
rect 29 703 279 750
rect 29 669 45 703
rect 263 669 279 703
rect 29 653 279 669
rect 337 703 587 750
rect 337 669 353 703
rect 571 669 587 703
rect 337 653 587 669
rect -587 585 -337 611
rect -279 585 -29 611
rect 29 585 279 611
rect 337 585 587 611
rect -587 -562 -337 -515
rect -587 -596 -571 -562
rect -353 -596 -337 -562
rect -587 -612 -337 -596
rect -279 -562 -29 -515
rect -279 -596 -263 -562
rect -45 -596 -29 -562
rect -279 -612 -29 -596
rect 29 -562 279 -515
rect 29 -596 45 -562
rect 263 -596 279 -562
rect 29 -612 279 -596
rect 337 -562 587 -515
rect 337 -596 353 -562
rect 571 -596 587 -562
rect 337 -612 587 -596
rect -587 -680 -337 -654
rect -279 -680 -29 -654
rect 29 -680 279 -654
rect 337 -680 587 -654
rect -587 -1827 -337 -1780
rect -587 -1861 -571 -1827
rect -353 -1861 -337 -1827
rect -587 -1877 -337 -1861
rect -279 -1827 -29 -1780
rect -279 -1861 -263 -1827
rect -45 -1861 -29 -1827
rect -279 -1877 -29 -1861
rect 29 -1827 279 -1780
rect 29 -1861 45 -1827
rect 263 -1861 279 -1827
rect 29 -1877 279 -1861
rect 337 -1827 587 -1780
rect 337 -1861 353 -1827
rect 571 -1861 587 -1827
rect 337 -1877 587 -1861
rect -587 -1945 -337 -1919
rect -279 -1945 -29 -1919
rect 29 -1945 279 -1919
rect 337 -1945 587 -1919
rect -587 -3092 -337 -3045
rect -587 -3126 -571 -3092
rect -353 -3126 -337 -3092
rect -587 -3142 -337 -3126
rect -279 -3092 -29 -3045
rect -279 -3126 -263 -3092
rect -45 -3126 -29 -3092
rect -279 -3142 -29 -3126
rect 29 -3092 279 -3045
rect 29 -3126 45 -3092
rect 263 -3126 279 -3092
rect 29 -3142 279 -3126
rect 337 -3092 587 -3045
rect 337 -3126 353 -3092
rect 571 -3126 587 -3092
rect 337 -3142 587 -3126
<< polycont >>
rect -571 1934 -353 1968
rect -263 1934 -45 1968
rect 45 1934 263 1968
rect 353 1934 571 1968
rect -571 669 -353 703
rect -263 669 -45 703
rect 45 669 263 703
rect 353 669 571 703
rect -571 -596 -353 -562
rect -263 -596 -45 -562
rect 45 -596 263 -562
rect 353 -596 571 -562
rect -571 -1861 -353 -1827
rect -263 -1861 -45 -1827
rect 45 -1861 263 -1827
rect 353 -1861 571 -1827
rect -571 -3126 -353 -3092
rect -263 -3126 -45 -3092
rect 45 -3126 263 -3092
rect 353 -3126 571 -3092
<< locali >>
rect -633 2834 -599 2850
rect -633 2280 -599 2296
rect -325 2834 -291 2850
rect -325 2280 -291 2296
rect -17 2834 17 2850
rect -17 2280 17 2296
rect 291 2834 325 2850
rect 291 2280 325 2296
rect 599 2834 633 2850
rect 599 2280 633 2296
rect -587 1934 -571 1968
rect -353 1934 -337 1968
rect -279 1934 -263 1968
rect -45 1934 -29 1968
rect 29 1934 45 1968
rect 263 1934 279 1968
rect 337 1934 353 1968
rect 571 1934 587 1968
rect -633 1569 -599 1585
rect -633 1015 -599 1031
rect -325 1569 -291 1585
rect -325 1015 -291 1031
rect -17 1569 17 1585
rect -17 1015 17 1031
rect 291 1569 325 1585
rect 291 1015 325 1031
rect 599 1569 633 1585
rect 599 1015 633 1031
rect -587 669 -571 703
rect -353 669 -337 703
rect -279 669 -263 703
rect -45 669 -29 703
rect 29 669 45 703
rect 263 669 279 703
rect 337 669 353 703
rect 571 669 587 703
rect -633 304 -599 320
rect -633 -250 -599 -234
rect -325 304 -291 320
rect -325 -250 -291 -234
rect -17 304 17 320
rect -17 -250 17 -234
rect 291 304 325 320
rect 291 -250 325 -234
rect 599 304 633 320
rect 599 -250 633 -234
rect -587 -596 -571 -562
rect -353 -596 -337 -562
rect -279 -596 -263 -562
rect -45 -596 -29 -562
rect 29 -596 45 -562
rect 263 -596 279 -562
rect 337 -596 353 -562
rect 571 -596 587 -562
rect -633 -961 -599 -945
rect -633 -1515 -599 -1499
rect -325 -961 -291 -945
rect -325 -1515 -291 -1499
rect -17 -961 17 -945
rect -17 -1515 17 -1499
rect 291 -961 325 -945
rect 291 -1515 325 -1499
rect 599 -961 633 -945
rect 599 -1515 633 -1499
rect -587 -1861 -571 -1827
rect -353 -1861 -337 -1827
rect -279 -1861 -263 -1827
rect -45 -1861 -29 -1827
rect 29 -1861 45 -1827
rect 263 -1861 279 -1827
rect 337 -1861 353 -1827
rect 571 -1861 587 -1827
rect -633 -2226 -599 -2210
rect -633 -2780 -599 -2764
rect -325 -2226 -291 -2210
rect -325 -2780 -291 -2764
rect -17 -2226 17 -2210
rect -17 -2780 17 -2764
rect 291 -2226 325 -2210
rect 291 -2780 325 -2764
rect 599 -2226 633 -2210
rect 599 -2780 633 -2764
rect -587 -3126 -571 -3092
rect -353 -3126 -337 -3092
rect -279 -3126 -263 -3092
rect -45 -3126 -29 -3092
rect 29 -3126 45 -3092
rect 263 -3126 279 -3092
rect 337 -3126 353 -3092
rect 571 -3126 587 -3092
<< viali >>
rect -633 2296 -599 2834
rect -325 2296 -291 2834
rect -17 2296 17 2834
rect 291 2296 325 2834
rect 599 2296 633 2834
rect -571 1934 -353 1968
rect -263 1934 -45 1968
rect 45 1934 263 1968
rect 353 1934 571 1968
rect -633 1031 -599 1569
rect -325 1031 -291 1569
rect -17 1031 17 1569
rect 291 1031 325 1569
rect 599 1031 633 1569
rect -571 669 -353 703
rect -263 669 -45 703
rect 45 669 263 703
rect 353 669 571 703
rect -633 -234 -599 304
rect -325 -234 -291 304
rect -17 -234 17 304
rect 291 -234 325 304
rect 599 -234 633 304
rect -571 -596 -353 -562
rect -263 -596 -45 -562
rect 45 -596 263 -562
rect 353 -596 571 -562
rect -633 -1499 -599 -961
rect -325 -1499 -291 -961
rect -17 -1499 17 -961
rect 291 -1499 325 -961
rect 599 -1499 633 -961
rect -571 -1861 -353 -1827
rect -263 -1861 -45 -1827
rect 45 -1861 263 -1827
rect 353 -1861 571 -1827
rect -633 -2764 -599 -2226
rect -325 -2764 -291 -2226
rect -17 -2764 17 -2226
rect 291 -2764 325 -2226
rect 599 -2764 633 -2226
rect -571 -3126 -353 -3092
rect -263 -3126 -45 -3092
rect 45 -3126 263 -3092
rect 353 -3126 571 -3092
<< metal1 >>
rect -639 2834 -593 2846
rect -639 2296 -633 2834
rect -599 2296 -593 2834
rect -639 2284 -593 2296
rect -331 2834 -285 2846
rect -331 2296 -325 2834
rect -291 2296 -285 2834
rect -331 2284 -285 2296
rect -23 2834 23 2846
rect -23 2296 -17 2834
rect 17 2296 23 2834
rect -23 2284 23 2296
rect 285 2834 331 2846
rect 285 2296 291 2834
rect 325 2296 331 2834
rect 285 2284 331 2296
rect 593 2834 639 2846
rect 593 2296 599 2834
rect 633 2296 639 2834
rect 593 2284 639 2296
rect -583 1968 -341 1974
rect -583 1934 -571 1968
rect -353 1934 -341 1968
rect -583 1928 -341 1934
rect -275 1968 -33 1974
rect -275 1934 -263 1968
rect -45 1934 -33 1968
rect -275 1928 -33 1934
rect 33 1968 275 1974
rect 33 1934 45 1968
rect 263 1934 275 1968
rect 33 1928 275 1934
rect 341 1968 583 1974
rect 341 1934 353 1968
rect 571 1934 583 1968
rect 341 1928 583 1934
rect -639 1569 -593 1581
rect -639 1031 -633 1569
rect -599 1031 -593 1569
rect -639 1019 -593 1031
rect -331 1569 -285 1581
rect -331 1031 -325 1569
rect -291 1031 -285 1569
rect -331 1019 -285 1031
rect -23 1569 23 1581
rect -23 1031 -17 1569
rect 17 1031 23 1569
rect -23 1019 23 1031
rect 285 1569 331 1581
rect 285 1031 291 1569
rect 325 1031 331 1569
rect 285 1019 331 1031
rect 593 1569 639 1581
rect 593 1031 599 1569
rect 633 1031 639 1569
rect 593 1019 639 1031
rect -583 703 -341 709
rect -583 669 -571 703
rect -353 669 -341 703
rect -583 663 -341 669
rect -275 703 -33 709
rect -275 669 -263 703
rect -45 669 -33 703
rect -275 663 -33 669
rect 33 703 275 709
rect 33 669 45 703
rect 263 669 275 703
rect 33 663 275 669
rect 341 703 583 709
rect 341 669 353 703
rect 571 669 583 703
rect 341 663 583 669
rect -639 304 -593 316
rect -639 -234 -633 304
rect -599 -234 -593 304
rect -639 -246 -593 -234
rect -331 304 -285 316
rect -331 -234 -325 304
rect -291 -234 -285 304
rect -331 -246 -285 -234
rect -23 304 23 316
rect -23 -234 -17 304
rect 17 -234 23 304
rect -23 -246 23 -234
rect 285 304 331 316
rect 285 -234 291 304
rect 325 -234 331 304
rect 285 -246 331 -234
rect 593 304 639 316
rect 593 -234 599 304
rect 633 -234 639 304
rect 593 -246 639 -234
rect -583 -562 -341 -556
rect -583 -596 -571 -562
rect -353 -596 -341 -562
rect -583 -602 -341 -596
rect -275 -562 -33 -556
rect -275 -596 -263 -562
rect -45 -596 -33 -562
rect -275 -602 -33 -596
rect 33 -562 275 -556
rect 33 -596 45 -562
rect 263 -596 275 -562
rect 33 -602 275 -596
rect 341 -562 583 -556
rect 341 -596 353 -562
rect 571 -596 583 -562
rect 341 -602 583 -596
rect -639 -961 -593 -949
rect -639 -1499 -633 -961
rect -599 -1499 -593 -961
rect -639 -1511 -593 -1499
rect -331 -961 -285 -949
rect -331 -1499 -325 -961
rect -291 -1499 -285 -961
rect -331 -1511 -285 -1499
rect -23 -961 23 -949
rect -23 -1499 -17 -961
rect 17 -1499 23 -961
rect -23 -1511 23 -1499
rect 285 -961 331 -949
rect 285 -1499 291 -961
rect 325 -1499 331 -961
rect 285 -1511 331 -1499
rect 593 -961 639 -949
rect 593 -1499 599 -961
rect 633 -1499 639 -961
rect 593 -1511 639 -1499
rect -583 -1827 -341 -1821
rect -583 -1861 -571 -1827
rect -353 -1861 -341 -1827
rect -583 -1867 -341 -1861
rect -275 -1827 -33 -1821
rect -275 -1861 -263 -1827
rect -45 -1861 -33 -1827
rect -275 -1867 -33 -1861
rect 33 -1827 275 -1821
rect 33 -1861 45 -1827
rect 263 -1861 275 -1827
rect 33 -1867 275 -1861
rect 341 -1827 583 -1821
rect 341 -1861 353 -1827
rect 571 -1861 583 -1827
rect 341 -1867 583 -1861
rect -639 -2226 -593 -2214
rect -639 -2764 -633 -2226
rect -599 -2764 -593 -2226
rect -639 -2776 -593 -2764
rect -331 -2226 -285 -2214
rect -331 -2764 -325 -2226
rect -291 -2764 -285 -2226
rect -331 -2776 -285 -2764
rect -23 -2226 23 -2214
rect -23 -2764 -17 -2226
rect 17 -2764 23 -2226
rect -23 -2776 23 -2764
rect 285 -2226 331 -2214
rect 285 -2764 291 -2226
rect 325 -2764 331 -2226
rect 285 -2776 331 -2764
rect 593 -2226 639 -2214
rect 593 -2764 599 -2226
rect 633 -2764 639 -2226
rect 593 -2776 639 -2764
rect -583 -3092 -341 -3086
rect -583 -3126 -571 -3092
rect -353 -3126 -341 -3092
rect -583 -3132 -341 -3126
rect -275 -3092 -33 -3086
rect -275 -3126 -263 -3092
rect -45 -3126 -33 -3092
rect -275 -3132 -33 -3126
rect 33 -3092 275 -3086
rect 33 -3126 45 -3092
rect 263 -3126 275 -3092
rect 33 -3132 275 -3126
rect 341 -3092 583 -3086
rect 341 -3126 353 -3092
rect 571 -3126 583 -3092
rect 341 -3132 583 -3126
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 5.5 l 1.25 m 5 nf 4 diffcov 50 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 class mosfet compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 50 viadrn 50 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1771413069
<< nwell >>
rect -5095 -563 5095 563
<< pmos >>
rect -4899 -344 -4649 344
rect -4591 -344 -4341 344
rect -4283 -344 -4033 344
rect -3975 -344 -3725 344
rect -3667 -344 -3417 344
rect -3359 -344 -3109 344
rect -3051 -344 -2801 344
rect -2743 -344 -2493 344
rect -2435 -344 -2185 344
rect -2127 -344 -1877 344
rect -1819 -344 -1569 344
rect -1511 -344 -1261 344
rect -1203 -344 -953 344
rect -895 -344 -645 344
rect -587 -344 -337 344
rect -279 -344 -29 344
rect 29 -344 279 344
rect 337 -344 587 344
rect 645 -344 895 344
rect 953 -344 1203 344
rect 1261 -344 1511 344
rect 1569 -344 1819 344
rect 1877 -344 2127 344
rect 2185 -344 2435 344
rect 2493 -344 2743 344
rect 2801 -344 3051 344
rect 3109 -344 3359 344
rect 3417 -344 3667 344
rect 3725 -344 3975 344
rect 4033 -344 4283 344
rect 4341 -344 4591 344
rect 4649 -344 4899 344
<< pdiff >>
rect -4957 332 -4899 344
rect -4957 -332 -4945 332
rect -4911 -332 -4899 332
rect -4957 -344 -4899 -332
rect -4649 332 -4591 344
rect -4649 -332 -4637 332
rect -4603 -332 -4591 332
rect -4649 -344 -4591 -332
rect -4341 332 -4283 344
rect -4341 -332 -4329 332
rect -4295 -332 -4283 332
rect -4341 -344 -4283 -332
rect -4033 332 -3975 344
rect -4033 -332 -4021 332
rect -3987 -332 -3975 332
rect -4033 -344 -3975 -332
rect -3725 332 -3667 344
rect -3725 -332 -3713 332
rect -3679 -332 -3667 332
rect -3725 -344 -3667 -332
rect -3417 332 -3359 344
rect -3417 -332 -3405 332
rect -3371 -332 -3359 332
rect -3417 -344 -3359 -332
rect -3109 332 -3051 344
rect -3109 -332 -3097 332
rect -3063 -332 -3051 332
rect -3109 -344 -3051 -332
rect -2801 332 -2743 344
rect -2801 -332 -2789 332
rect -2755 -332 -2743 332
rect -2801 -344 -2743 -332
rect -2493 332 -2435 344
rect -2493 -332 -2481 332
rect -2447 -332 -2435 332
rect -2493 -344 -2435 -332
rect -2185 332 -2127 344
rect -2185 -332 -2173 332
rect -2139 -332 -2127 332
rect -2185 -344 -2127 -332
rect -1877 332 -1819 344
rect -1877 -332 -1865 332
rect -1831 -332 -1819 332
rect -1877 -344 -1819 -332
rect -1569 332 -1511 344
rect -1569 -332 -1557 332
rect -1523 -332 -1511 332
rect -1569 -344 -1511 -332
rect -1261 332 -1203 344
rect -1261 -332 -1249 332
rect -1215 -332 -1203 332
rect -1261 -344 -1203 -332
rect -953 332 -895 344
rect -953 -332 -941 332
rect -907 -332 -895 332
rect -953 -344 -895 -332
rect -645 332 -587 344
rect -645 -332 -633 332
rect -599 -332 -587 332
rect -645 -344 -587 -332
rect -337 332 -279 344
rect -337 -332 -325 332
rect -291 -332 -279 332
rect -337 -344 -279 -332
rect -29 332 29 344
rect -29 -332 -17 332
rect 17 -332 29 332
rect -29 -344 29 -332
rect 279 332 337 344
rect 279 -332 291 332
rect 325 -332 337 332
rect 279 -344 337 -332
rect 587 332 645 344
rect 587 -332 599 332
rect 633 -332 645 332
rect 587 -344 645 -332
rect 895 332 953 344
rect 895 -332 907 332
rect 941 -332 953 332
rect 895 -344 953 -332
rect 1203 332 1261 344
rect 1203 -332 1215 332
rect 1249 -332 1261 332
rect 1203 -344 1261 -332
rect 1511 332 1569 344
rect 1511 -332 1523 332
rect 1557 -332 1569 332
rect 1511 -344 1569 -332
rect 1819 332 1877 344
rect 1819 -332 1831 332
rect 1865 -332 1877 332
rect 1819 -344 1877 -332
rect 2127 332 2185 344
rect 2127 -332 2139 332
rect 2173 -332 2185 332
rect 2127 -344 2185 -332
rect 2435 332 2493 344
rect 2435 -332 2447 332
rect 2481 -332 2493 332
rect 2435 -344 2493 -332
rect 2743 332 2801 344
rect 2743 -332 2755 332
rect 2789 -332 2801 332
rect 2743 -344 2801 -332
rect 3051 332 3109 344
rect 3051 -332 3063 332
rect 3097 -332 3109 332
rect 3051 -344 3109 -332
rect 3359 332 3417 344
rect 3359 -332 3371 332
rect 3405 -332 3417 332
rect 3359 -344 3417 -332
rect 3667 332 3725 344
rect 3667 -332 3679 332
rect 3713 -332 3725 332
rect 3667 -344 3725 -332
rect 3975 332 4033 344
rect 3975 -332 3987 332
rect 4021 -332 4033 332
rect 3975 -344 4033 -332
rect 4283 332 4341 344
rect 4283 -332 4295 332
rect 4329 -332 4341 332
rect 4283 -344 4341 -332
rect 4591 332 4649 344
rect 4591 -332 4603 332
rect 4637 -332 4649 332
rect 4591 -344 4649 -332
rect 4899 332 4957 344
rect 4899 -332 4911 332
rect 4945 -332 4957 332
rect 4899 -344 4957 -332
<< pdiffc >>
rect -4945 -332 -4911 332
rect -4637 -332 -4603 332
rect -4329 -332 -4295 332
rect -4021 -332 -3987 332
rect -3713 -332 -3679 332
rect -3405 -332 -3371 332
rect -3097 -332 -3063 332
rect -2789 -332 -2755 332
rect -2481 -332 -2447 332
rect -2173 -332 -2139 332
rect -1865 -332 -1831 332
rect -1557 -332 -1523 332
rect -1249 -332 -1215 332
rect -941 -332 -907 332
rect -633 -332 -599 332
rect -325 -332 -291 332
rect -17 -332 17 332
rect 291 -332 325 332
rect 599 -332 633 332
rect 907 -332 941 332
rect 1215 -332 1249 332
rect 1523 -332 1557 332
rect 1831 -332 1865 332
rect 2139 -332 2173 332
rect 2447 -332 2481 332
rect 2755 -332 2789 332
rect 3063 -332 3097 332
rect 3371 -332 3405 332
rect 3679 -332 3713 332
rect 3987 -332 4021 332
rect 4295 -332 4329 332
rect 4603 -332 4637 332
rect 4911 -332 4945 332
<< nsubdiff >>
rect -5059 493 -4963 527
rect 4963 493 5059 527
rect -5059 431 -5025 493
rect 5025 431 5059 493
rect -5059 -493 -5025 -431
rect 5025 -493 5059 -431
rect -5059 -527 -4963 -493
rect 4963 -527 5059 -493
<< nsubdiffcont >>
rect -4963 493 4963 527
rect -5059 -431 -5025 431
rect 5025 -431 5059 431
rect -4963 -527 4963 -493
<< poly >>
rect -4899 425 -4649 441
rect -4899 391 -4883 425
rect -4665 391 -4649 425
rect -4899 344 -4649 391
rect -4591 425 -4341 441
rect -4591 391 -4575 425
rect -4357 391 -4341 425
rect -4591 344 -4341 391
rect -4283 425 -4033 441
rect -4283 391 -4267 425
rect -4049 391 -4033 425
rect -4283 344 -4033 391
rect -3975 425 -3725 441
rect -3975 391 -3959 425
rect -3741 391 -3725 425
rect -3975 344 -3725 391
rect -3667 425 -3417 441
rect -3667 391 -3651 425
rect -3433 391 -3417 425
rect -3667 344 -3417 391
rect -3359 425 -3109 441
rect -3359 391 -3343 425
rect -3125 391 -3109 425
rect -3359 344 -3109 391
rect -3051 425 -2801 441
rect -3051 391 -3035 425
rect -2817 391 -2801 425
rect -3051 344 -2801 391
rect -2743 425 -2493 441
rect -2743 391 -2727 425
rect -2509 391 -2493 425
rect -2743 344 -2493 391
rect -2435 425 -2185 441
rect -2435 391 -2419 425
rect -2201 391 -2185 425
rect -2435 344 -2185 391
rect -2127 425 -1877 441
rect -2127 391 -2111 425
rect -1893 391 -1877 425
rect -2127 344 -1877 391
rect -1819 425 -1569 441
rect -1819 391 -1803 425
rect -1585 391 -1569 425
rect -1819 344 -1569 391
rect -1511 425 -1261 441
rect -1511 391 -1495 425
rect -1277 391 -1261 425
rect -1511 344 -1261 391
rect -1203 425 -953 441
rect -1203 391 -1187 425
rect -969 391 -953 425
rect -1203 344 -953 391
rect -895 425 -645 441
rect -895 391 -879 425
rect -661 391 -645 425
rect -895 344 -645 391
rect -587 425 -337 441
rect -587 391 -571 425
rect -353 391 -337 425
rect -587 344 -337 391
rect -279 425 -29 441
rect -279 391 -263 425
rect -45 391 -29 425
rect -279 344 -29 391
rect 29 425 279 441
rect 29 391 45 425
rect 263 391 279 425
rect 29 344 279 391
rect 337 425 587 441
rect 337 391 353 425
rect 571 391 587 425
rect 337 344 587 391
rect 645 425 895 441
rect 645 391 661 425
rect 879 391 895 425
rect 645 344 895 391
rect 953 425 1203 441
rect 953 391 969 425
rect 1187 391 1203 425
rect 953 344 1203 391
rect 1261 425 1511 441
rect 1261 391 1277 425
rect 1495 391 1511 425
rect 1261 344 1511 391
rect 1569 425 1819 441
rect 1569 391 1585 425
rect 1803 391 1819 425
rect 1569 344 1819 391
rect 1877 425 2127 441
rect 1877 391 1893 425
rect 2111 391 2127 425
rect 1877 344 2127 391
rect 2185 425 2435 441
rect 2185 391 2201 425
rect 2419 391 2435 425
rect 2185 344 2435 391
rect 2493 425 2743 441
rect 2493 391 2509 425
rect 2727 391 2743 425
rect 2493 344 2743 391
rect 2801 425 3051 441
rect 2801 391 2817 425
rect 3035 391 3051 425
rect 2801 344 3051 391
rect 3109 425 3359 441
rect 3109 391 3125 425
rect 3343 391 3359 425
rect 3109 344 3359 391
rect 3417 425 3667 441
rect 3417 391 3433 425
rect 3651 391 3667 425
rect 3417 344 3667 391
rect 3725 425 3975 441
rect 3725 391 3741 425
rect 3959 391 3975 425
rect 3725 344 3975 391
rect 4033 425 4283 441
rect 4033 391 4049 425
rect 4267 391 4283 425
rect 4033 344 4283 391
rect 4341 425 4591 441
rect 4341 391 4357 425
rect 4575 391 4591 425
rect 4341 344 4591 391
rect 4649 425 4899 441
rect 4649 391 4665 425
rect 4883 391 4899 425
rect 4649 344 4899 391
rect -4899 -391 -4649 -344
rect -4899 -425 -4883 -391
rect -4665 -425 -4649 -391
rect -4899 -441 -4649 -425
rect -4591 -391 -4341 -344
rect -4591 -425 -4575 -391
rect -4357 -425 -4341 -391
rect -4591 -441 -4341 -425
rect -4283 -391 -4033 -344
rect -4283 -425 -4267 -391
rect -4049 -425 -4033 -391
rect -4283 -441 -4033 -425
rect -3975 -391 -3725 -344
rect -3975 -425 -3959 -391
rect -3741 -425 -3725 -391
rect -3975 -441 -3725 -425
rect -3667 -391 -3417 -344
rect -3667 -425 -3651 -391
rect -3433 -425 -3417 -391
rect -3667 -441 -3417 -425
rect -3359 -391 -3109 -344
rect -3359 -425 -3343 -391
rect -3125 -425 -3109 -391
rect -3359 -441 -3109 -425
rect -3051 -391 -2801 -344
rect -3051 -425 -3035 -391
rect -2817 -425 -2801 -391
rect -3051 -441 -2801 -425
rect -2743 -391 -2493 -344
rect -2743 -425 -2727 -391
rect -2509 -425 -2493 -391
rect -2743 -441 -2493 -425
rect -2435 -391 -2185 -344
rect -2435 -425 -2419 -391
rect -2201 -425 -2185 -391
rect -2435 -441 -2185 -425
rect -2127 -391 -1877 -344
rect -2127 -425 -2111 -391
rect -1893 -425 -1877 -391
rect -2127 -441 -1877 -425
rect -1819 -391 -1569 -344
rect -1819 -425 -1803 -391
rect -1585 -425 -1569 -391
rect -1819 -441 -1569 -425
rect -1511 -391 -1261 -344
rect -1511 -425 -1495 -391
rect -1277 -425 -1261 -391
rect -1511 -441 -1261 -425
rect -1203 -391 -953 -344
rect -1203 -425 -1187 -391
rect -969 -425 -953 -391
rect -1203 -441 -953 -425
rect -895 -391 -645 -344
rect -895 -425 -879 -391
rect -661 -425 -645 -391
rect -895 -441 -645 -425
rect -587 -391 -337 -344
rect -587 -425 -571 -391
rect -353 -425 -337 -391
rect -587 -441 -337 -425
rect -279 -391 -29 -344
rect -279 -425 -263 -391
rect -45 -425 -29 -391
rect -279 -441 -29 -425
rect 29 -391 279 -344
rect 29 -425 45 -391
rect 263 -425 279 -391
rect 29 -441 279 -425
rect 337 -391 587 -344
rect 337 -425 353 -391
rect 571 -425 587 -391
rect 337 -441 587 -425
rect 645 -391 895 -344
rect 645 -425 661 -391
rect 879 -425 895 -391
rect 645 -441 895 -425
rect 953 -391 1203 -344
rect 953 -425 969 -391
rect 1187 -425 1203 -391
rect 953 -441 1203 -425
rect 1261 -391 1511 -344
rect 1261 -425 1277 -391
rect 1495 -425 1511 -391
rect 1261 -441 1511 -425
rect 1569 -391 1819 -344
rect 1569 -425 1585 -391
rect 1803 -425 1819 -391
rect 1569 -441 1819 -425
rect 1877 -391 2127 -344
rect 1877 -425 1893 -391
rect 2111 -425 2127 -391
rect 1877 -441 2127 -425
rect 2185 -391 2435 -344
rect 2185 -425 2201 -391
rect 2419 -425 2435 -391
rect 2185 -441 2435 -425
rect 2493 -391 2743 -344
rect 2493 -425 2509 -391
rect 2727 -425 2743 -391
rect 2493 -441 2743 -425
rect 2801 -391 3051 -344
rect 2801 -425 2817 -391
rect 3035 -425 3051 -391
rect 2801 -441 3051 -425
rect 3109 -391 3359 -344
rect 3109 -425 3125 -391
rect 3343 -425 3359 -391
rect 3109 -441 3359 -425
rect 3417 -391 3667 -344
rect 3417 -425 3433 -391
rect 3651 -425 3667 -391
rect 3417 -441 3667 -425
rect 3725 -391 3975 -344
rect 3725 -425 3741 -391
rect 3959 -425 3975 -391
rect 3725 -441 3975 -425
rect 4033 -391 4283 -344
rect 4033 -425 4049 -391
rect 4267 -425 4283 -391
rect 4033 -441 4283 -425
rect 4341 -391 4591 -344
rect 4341 -425 4357 -391
rect 4575 -425 4591 -391
rect 4341 -441 4591 -425
rect 4649 -391 4899 -344
rect 4649 -425 4665 -391
rect 4883 -425 4899 -391
rect 4649 -441 4899 -425
<< polycont >>
rect -4883 391 -4665 425
rect -4575 391 -4357 425
rect -4267 391 -4049 425
rect -3959 391 -3741 425
rect -3651 391 -3433 425
rect -3343 391 -3125 425
rect -3035 391 -2817 425
rect -2727 391 -2509 425
rect -2419 391 -2201 425
rect -2111 391 -1893 425
rect -1803 391 -1585 425
rect -1495 391 -1277 425
rect -1187 391 -969 425
rect -879 391 -661 425
rect -571 391 -353 425
rect -263 391 -45 425
rect 45 391 263 425
rect 353 391 571 425
rect 661 391 879 425
rect 969 391 1187 425
rect 1277 391 1495 425
rect 1585 391 1803 425
rect 1893 391 2111 425
rect 2201 391 2419 425
rect 2509 391 2727 425
rect 2817 391 3035 425
rect 3125 391 3343 425
rect 3433 391 3651 425
rect 3741 391 3959 425
rect 4049 391 4267 425
rect 4357 391 4575 425
rect 4665 391 4883 425
rect -4883 -425 -4665 -391
rect -4575 -425 -4357 -391
rect -4267 -425 -4049 -391
rect -3959 -425 -3741 -391
rect -3651 -425 -3433 -391
rect -3343 -425 -3125 -391
rect -3035 -425 -2817 -391
rect -2727 -425 -2509 -391
rect -2419 -425 -2201 -391
rect -2111 -425 -1893 -391
rect -1803 -425 -1585 -391
rect -1495 -425 -1277 -391
rect -1187 -425 -969 -391
rect -879 -425 -661 -391
rect -571 -425 -353 -391
rect -263 -425 -45 -391
rect 45 -425 263 -391
rect 353 -425 571 -391
rect 661 -425 879 -391
rect 969 -425 1187 -391
rect 1277 -425 1495 -391
rect 1585 -425 1803 -391
rect 1893 -425 2111 -391
rect 2201 -425 2419 -391
rect 2509 -425 2727 -391
rect 2817 -425 3035 -391
rect 3125 -425 3343 -391
rect 3433 -425 3651 -391
rect 3741 -425 3959 -391
rect 4049 -425 4267 -391
rect 4357 -425 4575 -391
rect 4665 -425 4883 -391
<< locali >>
rect -5059 493 -4963 527
rect 4963 493 5059 527
rect -5059 431 -5025 493
rect 5025 431 5059 493
rect -4899 391 -4883 425
rect -4665 391 -4649 425
rect -4591 391 -4575 425
rect -4357 391 -4341 425
rect -4283 391 -4267 425
rect -4049 391 -4033 425
rect -3975 391 -3959 425
rect -3741 391 -3725 425
rect -3667 391 -3651 425
rect -3433 391 -3417 425
rect -3359 391 -3343 425
rect -3125 391 -3109 425
rect -3051 391 -3035 425
rect -2817 391 -2801 425
rect -2743 391 -2727 425
rect -2509 391 -2493 425
rect -2435 391 -2419 425
rect -2201 391 -2185 425
rect -2127 391 -2111 425
rect -1893 391 -1877 425
rect -1819 391 -1803 425
rect -1585 391 -1569 425
rect -1511 391 -1495 425
rect -1277 391 -1261 425
rect -1203 391 -1187 425
rect -969 391 -953 425
rect -895 391 -879 425
rect -661 391 -645 425
rect -587 391 -571 425
rect -353 391 -337 425
rect -279 391 -263 425
rect -45 391 -29 425
rect 29 391 45 425
rect 263 391 279 425
rect 337 391 353 425
rect 571 391 587 425
rect 645 391 661 425
rect 879 391 895 425
rect 953 391 969 425
rect 1187 391 1203 425
rect 1261 391 1277 425
rect 1495 391 1511 425
rect 1569 391 1585 425
rect 1803 391 1819 425
rect 1877 391 1893 425
rect 2111 391 2127 425
rect 2185 391 2201 425
rect 2419 391 2435 425
rect 2493 391 2509 425
rect 2727 391 2743 425
rect 2801 391 2817 425
rect 3035 391 3051 425
rect 3109 391 3125 425
rect 3343 391 3359 425
rect 3417 391 3433 425
rect 3651 391 3667 425
rect 3725 391 3741 425
rect 3959 391 3975 425
rect 4033 391 4049 425
rect 4267 391 4283 425
rect 4341 391 4357 425
rect 4575 391 4591 425
rect 4649 391 4665 425
rect 4883 391 4899 425
rect -4945 332 -4911 348
rect -4945 -348 -4911 -332
rect -4637 332 -4603 348
rect -4637 -348 -4603 -332
rect -4329 332 -4295 348
rect -4329 -348 -4295 -332
rect -4021 332 -3987 348
rect -4021 -348 -3987 -332
rect -3713 332 -3679 348
rect -3713 -348 -3679 -332
rect -3405 332 -3371 348
rect -3405 -348 -3371 -332
rect -3097 332 -3063 348
rect -3097 -348 -3063 -332
rect -2789 332 -2755 348
rect -2789 -348 -2755 -332
rect -2481 332 -2447 348
rect -2481 -348 -2447 -332
rect -2173 332 -2139 348
rect -2173 -348 -2139 -332
rect -1865 332 -1831 348
rect -1865 -348 -1831 -332
rect -1557 332 -1523 348
rect -1557 -348 -1523 -332
rect -1249 332 -1215 348
rect -1249 -348 -1215 -332
rect -941 332 -907 348
rect -941 -348 -907 -332
rect -633 332 -599 348
rect -633 -348 -599 -332
rect -325 332 -291 348
rect -325 -348 -291 -332
rect -17 332 17 348
rect -17 -348 17 -332
rect 291 332 325 348
rect 291 -348 325 -332
rect 599 332 633 348
rect 599 -348 633 -332
rect 907 332 941 348
rect 907 -348 941 -332
rect 1215 332 1249 348
rect 1215 -348 1249 -332
rect 1523 332 1557 348
rect 1523 -348 1557 -332
rect 1831 332 1865 348
rect 1831 -348 1865 -332
rect 2139 332 2173 348
rect 2139 -348 2173 -332
rect 2447 332 2481 348
rect 2447 -348 2481 -332
rect 2755 332 2789 348
rect 2755 -348 2789 -332
rect 3063 332 3097 348
rect 3063 -348 3097 -332
rect 3371 332 3405 348
rect 3371 -348 3405 -332
rect 3679 332 3713 348
rect 3679 -348 3713 -332
rect 3987 332 4021 348
rect 3987 -348 4021 -332
rect 4295 332 4329 348
rect 4295 -348 4329 -332
rect 4603 332 4637 348
rect 4603 -348 4637 -332
rect 4911 332 4945 348
rect 4911 -348 4945 -332
rect -4899 -425 -4883 -391
rect -4665 -425 -4649 -391
rect -4591 -425 -4575 -391
rect -4357 -425 -4341 -391
rect -4283 -425 -4267 -391
rect -4049 -425 -4033 -391
rect -3975 -425 -3959 -391
rect -3741 -425 -3725 -391
rect -3667 -425 -3651 -391
rect -3433 -425 -3417 -391
rect -3359 -425 -3343 -391
rect -3125 -425 -3109 -391
rect -3051 -425 -3035 -391
rect -2817 -425 -2801 -391
rect -2743 -425 -2727 -391
rect -2509 -425 -2493 -391
rect -2435 -425 -2419 -391
rect -2201 -425 -2185 -391
rect -2127 -425 -2111 -391
rect -1893 -425 -1877 -391
rect -1819 -425 -1803 -391
rect -1585 -425 -1569 -391
rect -1511 -425 -1495 -391
rect -1277 -425 -1261 -391
rect -1203 -425 -1187 -391
rect -969 -425 -953 -391
rect -895 -425 -879 -391
rect -661 -425 -645 -391
rect -587 -425 -571 -391
rect -353 -425 -337 -391
rect -279 -425 -263 -391
rect -45 -425 -29 -391
rect 29 -425 45 -391
rect 263 -425 279 -391
rect 337 -425 353 -391
rect 571 -425 587 -391
rect 645 -425 661 -391
rect 879 -425 895 -391
rect 953 -425 969 -391
rect 1187 -425 1203 -391
rect 1261 -425 1277 -391
rect 1495 -425 1511 -391
rect 1569 -425 1585 -391
rect 1803 -425 1819 -391
rect 1877 -425 1893 -391
rect 2111 -425 2127 -391
rect 2185 -425 2201 -391
rect 2419 -425 2435 -391
rect 2493 -425 2509 -391
rect 2727 -425 2743 -391
rect 2801 -425 2817 -391
rect 3035 -425 3051 -391
rect 3109 -425 3125 -391
rect 3343 -425 3359 -391
rect 3417 -425 3433 -391
rect 3651 -425 3667 -391
rect 3725 -425 3741 -391
rect 3959 -425 3975 -391
rect 4033 -425 4049 -391
rect 4267 -425 4283 -391
rect 4341 -425 4357 -391
rect 4575 -425 4591 -391
rect 4649 -425 4665 -391
rect 4883 -425 4899 -391
rect -5059 -493 -5025 -431
rect 5025 -493 5059 -431
rect -5059 -527 -4963 -493
rect 4963 -527 5059 -493
<< viali >>
rect -4883 391 -4665 425
rect -4575 391 -4357 425
rect -4267 391 -4049 425
rect -3959 391 -3741 425
rect -3651 391 -3433 425
rect -3343 391 -3125 425
rect -3035 391 -2817 425
rect -2727 391 -2509 425
rect -2419 391 -2201 425
rect -2111 391 -1893 425
rect -1803 391 -1585 425
rect -1495 391 -1277 425
rect -1187 391 -969 425
rect -879 391 -661 425
rect -571 391 -353 425
rect -263 391 -45 425
rect 45 391 263 425
rect 353 391 571 425
rect 661 391 879 425
rect 969 391 1187 425
rect 1277 391 1495 425
rect 1585 391 1803 425
rect 1893 391 2111 425
rect 2201 391 2419 425
rect 2509 391 2727 425
rect 2817 391 3035 425
rect 3125 391 3343 425
rect 3433 391 3651 425
rect 3741 391 3959 425
rect 4049 391 4267 425
rect 4357 391 4575 425
rect 4665 391 4883 425
rect -4945 -332 -4911 332
rect -4637 -332 -4603 332
rect -4329 -332 -4295 332
rect -4021 -332 -3987 332
rect -3713 -332 -3679 332
rect -3405 -332 -3371 332
rect -3097 -332 -3063 332
rect -2789 -332 -2755 332
rect -2481 -332 -2447 332
rect -2173 -332 -2139 332
rect -1865 -332 -1831 332
rect -1557 -332 -1523 332
rect -1249 -332 -1215 332
rect -941 -332 -907 332
rect -633 -332 -599 332
rect -325 -332 -291 332
rect -17 -332 17 332
rect 291 -332 325 332
rect 599 -332 633 332
rect 907 -332 941 332
rect 1215 -332 1249 332
rect 1523 -332 1557 332
rect 1831 -332 1865 332
rect 2139 -332 2173 332
rect 2447 -332 2481 332
rect 2755 -332 2789 332
rect 3063 -332 3097 332
rect 3371 -332 3405 332
rect 3679 -332 3713 332
rect 3987 -332 4021 332
rect 4295 -332 4329 332
rect 4603 -332 4637 332
rect 4911 -332 4945 332
rect -4883 -425 -4665 -391
rect -4575 -425 -4357 -391
rect -4267 -425 -4049 -391
rect -3959 -425 -3741 -391
rect -3651 -425 -3433 -391
rect -3343 -425 -3125 -391
rect -3035 -425 -2817 -391
rect -2727 -425 -2509 -391
rect -2419 -425 -2201 -391
rect -2111 -425 -1893 -391
rect -1803 -425 -1585 -391
rect -1495 -425 -1277 -391
rect -1187 -425 -969 -391
rect -879 -425 -661 -391
rect -571 -425 -353 -391
rect -263 -425 -45 -391
rect 45 -425 263 -391
rect 353 -425 571 -391
rect 661 -425 879 -391
rect 969 -425 1187 -391
rect 1277 -425 1495 -391
rect 1585 -425 1803 -391
rect 1893 -425 2111 -391
rect 2201 -425 2419 -391
rect 2509 -425 2727 -391
rect 2817 -425 3035 -391
rect 3125 -425 3343 -391
rect 3433 -425 3651 -391
rect 3741 -425 3959 -391
rect 4049 -425 4267 -391
rect 4357 -425 4575 -391
rect 4665 -425 4883 -391
<< metal1 >>
rect -4895 425 -4653 431
rect -4895 391 -4883 425
rect -4665 391 -4653 425
rect -4895 385 -4653 391
rect -4587 425 -4345 431
rect -4587 391 -4575 425
rect -4357 391 -4345 425
rect -4587 385 -4345 391
rect -4279 425 -4037 431
rect -4279 391 -4267 425
rect -4049 391 -4037 425
rect -4279 385 -4037 391
rect -3971 425 -3729 431
rect -3971 391 -3959 425
rect -3741 391 -3729 425
rect -3971 385 -3729 391
rect -3663 425 -3421 431
rect -3663 391 -3651 425
rect -3433 391 -3421 425
rect -3663 385 -3421 391
rect -3355 425 -3113 431
rect -3355 391 -3343 425
rect -3125 391 -3113 425
rect -3355 385 -3113 391
rect -3047 425 -2805 431
rect -3047 391 -3035 425
rect -2817 391 -2805 425
rect -3047 385 -2805 391
rect -2739 425 -2497 431
rect -2739 391 -2727 425
rect -2509 391 -2497 425
rect -2739 385 -2497 391
rect -2431 425 -2189 431
rect -2431 391 -2419 425
rect -2201 391 -2189 425
rect -2431 385 -2189 391
rect -2123 425 -1881 431
rect -2123 391 -2111 425
rect -1893 391 -1881 425
rect -2123 385 -1881 391
rect -1815 425 -1573 431
rect -1815 391 -1803 425
rect -1585 391 -1573 425
rect -1815 385 -1573 391
rect -1507 425 -1265 431
rect -1507 391 -1495 425
rect -1277 391 -1265 425
rect -1507 385 -1265 391
rect -1199 425 -957 431
rect -1199 391 -1187 425
rect -969 391 -957 425
rect -1199 385 -957 391
rect -891 425 -649 431
rect -891 391 -879 425
rect -661 391 -649 425
rect -891 385 -649 391
rect -583 425 -341 431
rect -583 391 -571 425
rect -353 391 -341 425
rect -583 385 -341 391
rect -275 425 -33 431
rect -275 391 -263 425
rect -45 391 -33 425
rect -275 385 -33 391
rect 33 425 275 431
rect 33 391 45 425
rect 263 391 275 425
rect 33 385 275 391
rect 341 425 583 431
rect 341 391 353 425
rect 571 391 583 425
rect 341 385 583 391
rect 649 425 891 431
rect 649 391 661 425
rect 879 391 891 425
rect 649 385 891 391
rect 957 425 1199 431
rect 957 391 969 425
rect 1187 391 1199 425
rect 957 385 1199 391
rect 1265 425 1507 431
rect 1265 391 1277 425
rect 1495 391 1507 425
rect 1265 385 1507 391
rect 1573 425 1815 431
rect 1573 391 1585 425
rect 1803 391 1815 425
rect 1573 385 1815 391
rect 1881 425 2123 431
rect 1881 391 1893 425
rect 2111 391 2123 425
rect 1881 385 2123 391
rect 2189 425 2431 431
rect 2189 391 2201 425
rect 2419 391 2431 425
rect 2189 385 2431 391
rect 2497 425 2739 431
rect 2497 391 2509 425
rect 2727 391 2739 425
rect 2497 385 2739 391
rect 2805 425 3047 431
rect 2805 391 2817 425
rect 3035 391 3047 425
rect 2805 385 3047 391
rect 3113 425 3355 431
rect 3113 391 3125 425
rect 3343 391 3355 425
rect 3113 385 3355 391
rect 3421 425 3663 431
rect 3421 391 3433 425
rect 3651 391 3663 425
rect 3421 385 3663 391
rect 3729 425 3971 431
rect 3729 391 3741 425
rect 3959 391 3971 425
rect 3729 385 3971 391
rect 4037 425 4279 431
rect 4037 391 4049 425
rect 4267 391 4279 425
rect 4037 385 4279 391
rect 4345 425 4587 431
rect 4345 391 4357 425
rect 4575 391 4587 425
rect 4345 385 4587 391
rect 4653 425 4895 431
rect 4653 391 4665 425
rect 4883 391 4895 425
rect 4653 385 4895 391
rect -4951 332 -4905 344
rect -4951 -332 -4945 332
rect -4911 -332 -4905 332
rect -4951 -344 -4905 -332
rect -4643 332 -4597 344
rect -4643 -332 -4637 332
rect -4603 -332 -4597 332
rect -4643 -344 -4597 -332
rect -4335 332 -4289 344
rect -4335 -332 -4329 332
rect -4295 -332 -4289 332
rect -4335 -344 -4289 -332
rect -4027 332 -3981 344
rect -4027 -332 -4021 332
rect -3987 -332 -3981 332
rect -4027 -344 -3981 -332
rect -3719 332 -3673 344
rect -3719 -332 -3713 332
rect -3679 -332 -3673 332
rect -3719 -344 -3673 -332
rect -3411 332 -3365 344
rect -3411 -332 -3405 332
rect -3371 -332 -3365 332
rect -3411 -344 -3365 -332
rect -3103 332 -3057 344
rect -3103 -332 -3097 332
rect -3063 -332 -3057 332
rect -3103 -344 -3057 -332
rect -2795 332 -2749 344
rect -2795 -332 -2789 332
rect -2755 -332 -2749 332
rect -2795 -344 -2749 -332
rect -2487 332 -2441 344
rect -2487 -332 -2481 332
rect -2447 -332 -2441 332
rect -2487 -344 -2441 -332
rect -2179 332 -2133 344
rect -2179 -332 -2173 332
rect -2139 -332 -2133 332
rect -2179 -344 -2133 -332
rect -1871 332 -1825 344
rect -1871 -332 -1865 332
rect -1831 -332 -1825 332
rect -1871 -344 -1825 -332
rect -1563 332 -1517 344
rect -1563 -332 -1557 332
rect -1523 -332 -1517 332
rect -1563 -344 -1517 -332
rect -1255 332 -1209 344
rect -1255 -332 -1249 332
rect -1215 -332 -1209 332
rect -1255 -344 -1209 -332
rect -947 332 -901 344
rect -947 -332 -941 332
rect -907 -332 -901 332
rect -947 -344 -901 -332
rect -639 332 -593 344
rect -639 -332 -633 332
rect -599 -332 -593 332
rect -639 -344 -593 -332
rect -331 332 -285 344
rect -331 -332 -325 332
rect -291 -332 -285 332
rect -331 -344 -285 -332
rect -23 332 23 344
rect -23 -332 -17 332
rect 17 -332 23 332
rect -23 -344 23 -332
rect 285 332 331 344
rect 285 -332 291 332
rect 325 -332 331 332
rect 285 -344 331 -332
rect 593 332 639 344
rect 593 -332 599 332
rect 633 -332 639 332
rect 593 -344 639 -332
rect 901 332 947 344
rect 901 -332 907 332
rect 941 -332 947 332
rect 901 -344 947 -332
rect 1209 332 1255 344
rect 1209 -332 1215 332
rect 1249 -332 1255 332
rect 1209 -344 1255 -332
rect 1517 332 1563 344
rect 1517 -332 1523 332
rect 1557 -332 1563 332
rect 1517 -344 1563 -332
rect 1825 332 1871 344
rect 1825 -332 1831 332
rect 1865 -332 1871 332
rect 1825 -344 1871 -332
rect 2133 332 2179 344
rect 2133 -332 2139 332
rect 2173 -332 2179 332
rect 2133 -344 2179 -332
rect 2441 332 2487 344
rect 2441 -332 2447 332
rect 2481 -332 2487 332
rect 2441 -344 2487 -332
rect 2749 332 2795 344
rect 2749 -332 2755 332
rect 2789 -332 2795 332
rect 2749 -344 2795 -332
rect 3057 332 3103 344
rect 3057 -332 3063 332
rect 3097 -332 3103 332
rect 3057 -344 3103 -332
rect 3365 332 3411 344
rect 3365 -332 3371 332
rect 3405 -332 3411 332
rect 3365 -344 3411 -332
rect 3673 332 3719 344
rect 3673 -332 3679 332
rect 3713 -332 3719 332
rect 3673 -344 3719 -332
rect 3981 332 4027 344
rect 3981 -332 3987 332
rect 4021 -332 4027 332
rect 3981 -344 4027 -332
rect 4289 332 4335 344
rect 4289 -332 4295 332
rect 4329 -332 4335 332
rect 4289 -344 4335 -332
rect 4597 332 4643 344
rect 4597 -332 4603 332
rect 4637 -332 4643 332
rect 4597 -344 4643 -332
rect 4905 332 4951 344
rect 4905 -332 4911 332
rect 4945 -332 4951 332
rect 4905 -344 4951 -332
rect -4895 -391 -4653 -385
rect -4895 -425 -4883 -391
rect -4665 -425 -4653 -391
rect -4895 -431 -4653 -425
rect -4587 -391 -4345 -385
rect -4587 -425 -4575 -391
rect -4357 -425 -4345 -391
rect -4587 -431 -4345 -425
rect -4279 -391 -4037 -385
rect -4279 -425 -4267 -391
rect -4049 -425 -4037 -391
rect -4279 -431 -4037 -425
rect -3971 -391 -3729 -385
rect -3971 -425 -3959 -391
rect -3741 -425 -3729 -391
rect -3971 -431 -3729 -425
rect -3663 -391 -3421 -385
rect -3663 -425 -3651 -391
rect -3433 -425 -3421 -391
rect -3663 -431 -3421 -425
rect -3355 -391 -3113 -385
rect -3355 -425 -3343 -391
rect -3125 -425 -3113 -391
rect -3355 -431 -3113 -425
rect -3047 -391 -2805 -385
rect -3047 -425 -3035 -391
rect -2817 -425 -2805 -391
rect -3047 -431 -2805 -425
rect -2739 -391 -2497 -385
rect -2739 -425 -2727 -391
rect -2509 -425 -2497 -391
rect -2739 -431 -2497 -425
rect -2431 -391 -2189 -385
rect -2431 -425 -2419 -391
rect -2201 -425 -2189 -391
rect -2431 -431 -2189 -425
rect -2123 -391 -1881 -385
rect -2123 -425 -2111 -391
rect -1893 -425 -1881 -391
rect -2123 -431 -1881 -425
rect -1815 -391 -1573 -385
rect -1815 -425 -1803 -391
rect -1585 -425 -1573 -391
rect -1815 -431 -1573 -425
rect -1507 -391 -1265 -385
rect -1507 -425 -1495 -391
rect -1277 -425 -1265 -391
rect -1507 -431 -1265 -425
rect -1199 -391 -957 -385
rect -1199 -425 -1187 -391
rect -969 -425 -957 -391
rect -1199 -431 -957 -425
rect -891 -391 -649 -385
rect -891 -425 -879 -391
rect -661 -425 -649 -391
rect -891 -431 -649 -425
rect -583 -391 -341 -385
rect -583 -425 -571 -391
rect -353 -425 -341 -391
rect -583 -431 -341 -425
rect -275 -391 -33 -385
rect -275 -425 -263 -391
rect -45 -425 -33 -391
rect -275 -431 -33 -425
rect 33 -391 275 -385
rect 33 -425 45 -391
rect 263 -425 275 -391
rect 33 -431 275 -425
rect 341 -391 583 -385
rect 341 -425 353 -391
rect 571 -425 583 -391
rect 341 -431 583 -425
rect 649 -391 891 -385
rect 649 -425 661 -391
rect 879 -425 891 -391
rect 649 -431 891 -425
rect 957 -391 1199 -385
rect 957 -425 969 -391
rect 1187 -425 1199 -391
rect 957 -431 1199 -425
rect 1265 -391 1507 -385
rect 1265 -425 1277 -391
rect 1495 -425 1507 -391
rect 1265 -431 1507 -425
rect 1573 -391 1815 -385
rect 1573 -425 1585 -391
rect 1803 -425 1815 -391
rect 1573 -431 1815 -425
rect 1881 -391 2123 -385
rect 1881 -425 1893 -391
rect 2111 -425 2123 -391
rect 1881 -431 2123 -425
rect 2189 -391 2431 -385
rect 2189 -425 2201 -391
rect 2419 -425 2431 -391
rect 2189 -431 2431 -425
rect 2497 -391 2739 -385
rect 2497 -425 2509 -391
rect 2727 -425 2739 -391
rect 2497 -431 2739 -425
rect 2805 -391 3047 -385
rect 2805 -425 2817 -391
rect 3035 -425 3047 -391
rect 2805 -431 3047 -425
rect 3113 -391 3355 -385
rect 3113 -425 3125 -391
rect 3343 -425 3355 -391
rect 3113 -431 3355 -425
rect 3421 -391 3663 -385
rect 3421 -425 3433 -391
rect 3651 -425 3663 -391
rect 3421 -431 3663 -425
rect 3729 -391 3971 -385
rect 3729 -425 3741 -391
rect 3959 -425 3971 -391
rect 3729 -431 3971 -425
rect 4037 -391 4279 -385
rect 4037 -425 4049 -391
rect 4267 -425 4279 -391
rect 4037 -431 4279 -425
rect 4345 -391 4587 -385
rect 4345 -425 4357 -391
rect 4575 -425 4587 -391
rect 4345 -431 4587 -425
rect 4653 -391 4895 -385
rect 4653 -425 4665 -391
rect 4883 -425 4895 -391
rect 4653 -431 4895 -425
<< properties >>
string FIXED_BBOX -5042 -510 5042 510
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 3.4375 l 1.25 m 1 nf 32 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 class mosfet compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1770979109
<< nwell >>
rect -4297 -564 4297 598
<< pmos >>
rect -4203 -464 -3203 536
rect -3145 -464 -2145 536
rect -2087 -464 -1087 536
rect -1029 -464 -29 536
rect 29 -464 1029 536
rect 1087 -464 2087 536
rect 2145 -464 3145 536
rect 3203 -464 4203 536
<< pdiff >>
rect -4261 524 -4203 536
rect -4261 -452 -4249 524
rect -4215 -452 -4203 524
rect -4261 -464 -4203 -452
rect -3203 524 -3145 536
rect -3203 -452 -3191 524
rect -3157 -452 -3145 524
rect -3203 -464 -3145 -452
rect -2145 524 -2087 536
rect -2145 -452 -2133 524
rect -2099 -452 -2087 524
rect -2145 -464 -2087 -452
rect -1087 524 -1029 536
rect -1087 -452 -1075 524
rect -1041 -452 -1029 524
rect -1087 -464 -1029 -452
rect -29 524 29 536
rect -29 -452 -17 524
rect 17 -452 29 524
rect -29 -464 29 -452
rect 1029 524 1087 536
rect 1029 -452 1041 524
rect 1075 -452 1087 524
rect 1029 -464 1087 -452
rect 2087 524 2145 536
rect 2087 -452 2099 524
rect 2133 -452 2145 524
rect 2087 -464 2145 -452
rect 3145 524 3203 536
rect 3145 -452 3157 524
rect 3191 -452 3203 524
rect 3145 -464 3203 -452
rect 4203 524 4261 536
rect 4203 -452 4215 524
rect 4249 -452 4261 524
rect 4203 -464 4261 -452
<< pdiffc >>
rect -4249 -452 -4215 524
rect -3191 -452 -3157 524
rect -2133 -452 -2099 524
rect -1075 -452 -1041 524
rect -17 -452 17 524
rect 1041 -452 1075 524
rect 2099 -452 2133 524
rect 3157 -452 3191 524
rect 4215 -452 4249 524
<< poly >>
rect -4203 536 -3203 562
rect -3145 536 -2145 562
rect -2087 536 -1087 562
rect -1029 536 -29 562
rect 29 536 1029 562
rect 1087 536 2087 562
rect 2145 536 3145 562
rect 3203 536 4203 562
rect -4203 -511 -3203 -464
rect -4203 -545 -4187 -511
rect -3219 -545 -3203 -511
rect -4203 -561 -3203 -545
rect -3145 -511 -2145 -464
rect -3145 -545 -3129 -511
rect -2161 -545 -2145 -511
rect -3145 -561 -2145 -545
rect -2087 -511 -1087 -464
rect -2087 -545 -2071 -511
rect -1103 -545 -1087 -511
rect -2087 -561 -1087 -545
rect -1029 -511 -29 -464
rect -1029 -545 -1013 -511
rect -45 -545 -29 -511
rect -1029 -561 -29 -545
rect 29 -511 1029 -464
rect 29 -545 45 -511
rect 1013 -545 1029 -511
rect 29 -561 1029 -545
rect 1087 -511 2087 -464
rect 1087 -545 1103 -511
rect 2071 -545 2087 -511
rect 1087 -561 2087 -545
rect 2145 -511 3145 -464
rect 2145 -545 2161 -511
rect 3129 -545 3145 -511
rect 2145 -561 3145 -545
rect 3203 -511 4203 -464
rect 3203 -545 3219 -511
rect 4187 -545 4203 -511
rect 3203 -561 4203 -545
<< polycont >>
rect -4187 -545 -3219 -511
rect -3129 -545 -2161 -511
rect -2071 -545 -1103 -511
rect -1013 -545 -45 -511
rect 45 -545 1013 -511
rect 1103 -545 2071 -511
rect 2161 -545 3129 -511
rect 3219 -545 4187 -511
<< locali >>
rect -4249 524 -4215 540
rect -4249 -468 -4215 -452
rect -3191 524 -3157 540
rect -3191 -468 -3157 -452
rect -2133 524 -2099 540
rect -2133 -468 -2099 -452
rect -1075 524 -1041 540
rect -1075 -468 -1041 -452
rect -17 524 17 540
rect -17 -468 17 -452
rect 1041 524 1075 540
rect 1041 -468 1075 -452
rect 2099 524 2133 540
rect 2099 -468 2133 -452
rect 3157 524 3191 540
rect 3157 -468 3191 -452
rect 4215 524 4249 540
rect 4215 -468 4249 -452
rect -4203 -545 -4187 -511
rect -3219 -545 -3203 -511
rect -3145 -545 -3129 -511
rect -2161 -545 -2145 -511
rect -2087 -545 -2071 -511
rect -1103 -545 -1087 -511
rect -1029 -545 -1013 -511
rect -45 -545 -29 -511
rect 29 -545 45 -511
rect 1013 -545 1029 -511
rect 1087 -545 1103 -511
rect 2071 -545 2087 -511
rect 2145 -545 2161 -511
rect 3129 -545 3145 -511
rect 3203 -545 3219 -511
rect 4187 -545 4203 -511
<< viali >>
rect -4249 -452 -4215 524
rect -3191 -452 -3157 524
rect -2133 -452 -2099 524
rect -1075 -452 -1041 524
rect -17 -452 17 524
rect 1041 -452 1075 524
rect 2099 -452 2133 524
rect 3157 -452 3191 524
rect 4215 -452 4249 524
rect -4187 -545 -3219 -511
rect -3129 -545 -2161 -511
rect -2071 -545 -1103 -511
rect -1013 -545 -45 -511
rect 45 -545 1013 -511
rect 1103 -545 2071 -511
rect 2161 -545 3129 -511
rect 3219 -545 4187 -511
<< metal1 >>
rect -4255 524 -4209 536
rect -4255 -452 -4249 524
rect -4215 -452 -4209 524
rect -4255 -464 -4209 -452
rect -3197 524 -3151 536
rect -3197 -452 -3191 524
rect -3157 -452 -3151 524
rect -3197 -464 -3151 -452
rect -2139 524 -2093 536
rect -2139 -452 -2133 524
rect -2099 -452 -2093 524
rect -2139 -464 -2093 -452
rect -1081 524 -1035 536
rect -1081 -452 -1075 524
rect -1041 -452 -1035 524
rect -1081 -464 -1035 -452
rect -23 524 23 536
rect -23 -452 -17 524
rect 17 -452 23 524
rect -23 -464 23 -452
rect 1035 524 1081 536
rect 1035 -452 1041 524
rect 1075 -452 1081 524
rect 1035 -464 1081 -452
rect 2093 524 2139 536
rect 2093 -452 2099 524
rect 2133 -452 2139 524
rect 2093 -464 2139 -452
rect 3151 524 3197 536
rect 3151 -452 3157 524
rect 3191 -452 3197 524
rect 3151 -464 3197 -452
rect 4209 524 4255 536
rect 4209 -452 4215 524
rect 4249 -452 4255 524
rect 4209 -464 4255 -452
rect -4199 -511 -3207 -505
rect -4199 -545 -4187 -511
rect -3219 -545 -3207 -511
rect -4199 -551 -3207 -545
rect -3141 -511 -2149 -505
rect -3141 -545 -3129 -511
rect -2161 -545 -2149 -511
rect -3141 -551 -2149 -545
rect -2083 -511 -1091 -505
rect -2083 -545 -2071 -511
rect -1103 -545 -1091 -511
rect -2083 -551 -1091 -545
rect -1025 -511 -33 -505
rect -1025 -545 -1013 -511
rect -45 -545 -33 -511
rect -1025 -551 -33 -545
rect 33 -511 1025 -505
rect 33 -545 45 -511
rect 1013 -545 1025 -511
rect 33 -551 1025 -545
rect 1091 -511 2083 -505
rect 1091 -545 1103 -511
rect 2071 -545 2083 -511
rect 1091 -551 2083 -545
rect 2149 -511 3141 -505
rect 2149 -545 2161 -511
rect 3129 -545 3141 -511
rect 2149 -551 3141 -545
rect 3207 -511 4199 -505
rect 3207 -545 3219 -511
rect 4187 -545 4199 -511
rect 3207 -551 4199 -545
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 5.0 l 5.0 m 1 nf 8 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 class mosfet compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1771414049
<< metal3 >>
rect -3492 1512 -120 1540
rect -3492 -1512 -204 1512
rect -140 -1512 -120 1512
rect -3492 -1540 -120 -1512
rect 120 1512 3492 1540
rect 120 -1512 3408 1512
rect 3472 -1512 3492 1512
rect 120 -1540 3492 -1512
<< via3 >>
rect -204 -1512 -140 1512
rect 3408 -1512 3472 1512
<< mimcap >>
rect -3452 1460 -452 1500
rect -3452 -1460 -3412 1460
rect -492 -1460 -452 1460
rect -3452 -1500 -452 -1460
rect 160 1460 3160 1500
rect 160 -1460 200 1460
rect 3120 -1460 3160 1460
rect 160 -1500 3160 -1460
<< mimcapcontact >>
rect -3412 -1460 -492 1460
rect 200 -1460 3120 1460
<< metal4 >>
rect -220 1512 -124 1528
rect -3413 1460 -491 1461
rect -3413 -1460 -3412 1460
rect -492 -1460 -491 1460
rect -3413 -1461 -491 -1460
rect -220 -1512 -204 1512
rect -140 -1512 -124 1512
rect 3392 1512 3488 1528
rect 199 1460 3121 1461
rect 199 -1460 200 1460
rect 3120 -1460 3121 1460
rect 199 -1461 3121 -1460
rect -220 -1528 -124 -1512
rect 3392 -1512 3408 1512
rect 3472 -1512 3488 1512
rect 3392 -1528 3488 -1512
<< properties >>
string FIXED_BBOX 120 -1540 3200 1540
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 15.0 l 15.0 val 461.4 carea 2.00 cperi 0.19 class capacitor nx 2 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>

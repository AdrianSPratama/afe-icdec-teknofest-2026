magic
tech sky130A
magscale 1 2
timestamp 1771116256
<< pwell >>
rect -783 -510 783 510
<< nmos >>
rect -587 -300 -337 300
rect -279 -300 -29 300
rect 29 -300 279 300
rect 337 -300 587 300
<< ndiff >>
rect -645 288 -587 300
rect -645 -288 -633 288
rect -599 -288 -587 288
rect -645 -300 -587 -288
rect -337 288 -279 300
rect -337 -288 -325 288
rect -291 -288 -279 288
rect -337 -300 -279 -288
rect -29 288 29 300
rect -29 -288 -17 288
rect 17 -288 29 288
rect -29 -300 29 -288
rect 279 288 337 300
rect 279 -288 291 288
rect 325 -288 337 288
rect 279 -300 337 -288
rect 587 288 645 300
rect 587 -288 599 288
rect 633 -288 645 288
rect 587 -300 645 -288
<< ndiffc >>
rect -633 -288 -599 288
rect -325 -288 -291 288
rect -17 -288 17 288
rect 291 -288 325 288
rect 599 -288 633 288
<< psubdiff >>
rect -747 440 -651 474
rect 651 440 747 474
rect -747 378 -713 440
rect 713 378 747 440
rect -747 -440 -713 -378
rect 713 -440 747 -378
rect -747 -474 -651 -440
rect 651 -474 747 -440
<< psubdiffcont >>
rect -651 440 651 474
rect -747 -378 -713 378
rect 713 -378 747 378
rect -651 -474 651 -440
<< poly >>
rect -587 372 -337 388
rect -587 338 -571 372
rect -353 338 -337 372
rect -587 300 -337 338
rect -279 372 -29 388
rect -279 338 -263 372
rect -45 338 -29 372
rect -279 300 -29 338
rect 29 372 279 388
rect 29 338 45 372
rect 263 338 279 372
rect 29 300 279 338
rect 337 372 587 388
rect 337 338 353 372
rect 571 338 587 372
rect 337 300 587 338
rect -587 -338 -337 -300
rect -587 -372 -571 -338
rect -353 -372 -337 -338
rect -587 -388 -337 -372
rect -279 -338 -29 -300
rect -279 -372 -263 -338
rect -45 -372 -29 -338
rect -279 -388 -29 -372
rect 29 -338 279 -300
rect 29 -372 45 -338
rect 263 -372 279 -338
rect 29 -388 279 -372
rect 337 -338 587 -300
rect 337 -372 353 -338
rect 571 -372 587 -338
rect 337 -388 587 -372
<< polycont >>
rect -571 338 -353 372
rect -263 338 -45 372
rect 45 338 263 372
rect 353 338 571 372
rect -571 -372 -353 -338
rect -263 -372 -45 -338
rect 45 -372 263 -338
rect 353 -372 571 -338
<< locali >>
rect -747 440 -651 474
rect 651 440 747 474
rect -747 378 -713 440
rect 713 378 747 440
rect -587 338 -571 372
rect -353 338 -337 372
rect -279 338 -263 372
rect -45 338 -29 372
rect 29 338 45 372
rect 263 338 279 372
rect 337 338 353 372
rect 571 338 587 372
rect -633 288 -599 304
rect -633 -304 -599 -288
rect -325 288 -291 304
rect -325 -304 -291 -288
rect -17 288 17 304
rect -17 -304 17 -288
rect 291 288 325 304
rect 291 -304 325 -288
rect 599 288 633 304
rect 599 -304 633 -288
rect -587 -372 -571 -338
rect -353 -372 -337 -338
rect -279 -372 -263 -338
rect -45 -372 -29 -338
rect 29 -372 45 -338
rect 263 -372 279 -338
rect 337 -372 353 -338
rect 571 -372 587 -338
rect -747 -440 -713 -378
rect 713 -440 747 -378
rect -747 -474 -651 -440
rect 651 -474 747 -440
<< viali >>
rect -571 338 -353 372
rect -263 338 -45 372
rect 45 338 263 372
rect 353 338 571 372
rect -633 -288 -599 288
rect -325 -288 -291 288
rect -17 -288 17 288
rect 291 -288 325 288
rect 599 -288 633 288
rect -571 -372 -353 -338
rect -263 -372 -45 -338
rect 45 -372 263 -338
rect 353 -372 571 -338
<< metal1 >>
rect -583 372 -341 378
rect -583 338 -571 372
rect -353 338 -341 372
rect -583 332 -341 338
rect -275 372 -33 378
rect -275 338 -263 372
rect -45 338 -33 372
rect -275 332 -33 338
rect 33 372 275 378
rect 33 338 45 372
rect 263 338 275 372
rect 33 332 275 338
rect 341 372 583 378
rect 341 338 353 372
rect 571 338 583 372
rect 341 332 583 338
rect -639 288 -593 300
rect -639 -288 -633 288
rect -599 -288 -593 288
rect -639 -300 -593 -288
rect -331 288 -285 300
rect -331 -288 -325 288
rect -291 -288 -285 288
rect -331 -300 -285 -288
rect -23 288 23 300
rect -23 -288 -17 288
rect 17 -288 23 288
rect -23 -300 23 -288
rect 285 288 331 300
rect 285 -288 291 288
rect 325 -288 331 288
rect 285 -300 331 -288
rect 593 288 639 300
rect 593 -288 599 288
rect 633 -288 639 288
rect 593 -300 639 -288
rect -583 -338 -341 -332
rect -583 -372 -571 -338
rect -353 -372 -341 -338
rect -583 -378 -341 -372
rect -275 -338 -33 -332
rect -275 -372 -263 -338
rect -45 -372 -33 -338
rect -275 -378 -33 -372
rect 33 -338 275 -332
rect 33 -372 45 -338
rect 263 -372 275 -338
rect 33 -378 275 -372
rect 341 -338 583 -332
rect 341 -372 353 -338
rect 571 -372 583 -338
rect 341 -378 583 -372
<< properties >>
string FIXED_BBOX -730 -457 730 457
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 3.0 l 1.25 m 1 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 class mosfet compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

magic
tech sky130A
magscale 1 10
timestamp 1771420802
<< error_p >>
rect -4590 16520 4590 16580
rect -4590 -16520 -4530 16520
rect -4410 16340 4410 16400
rect -4410 15820 -4350 16340
rect -4345 15820 -4265 15900
rect -4195 15820 -4115 15900
rect 4115 15820 4195 15900
rect 4265 15820 4345 15900
rect 4350 15820 4410 16340
rect -4425 15740 -4345 15820
rect -4115 15740 -4035 15820
rect 4035 15740 4115 15820
rect 4345 15740 4425 15820
rect -4410 -15740 -4350 15740
rect -3655 14302 -3575 14382
rect -3505 14302 -3425 14382
rect -1885 14302 -1805 14382
rect -1735 14302 -1655 14382
rect -115 14302 -35 14382
rect 35 14302 115 14382
rect 1655 14302 1735 14382
rect 1805 14302 1885 14382
rect 3425 14302 3505 14382
rect 3575 14302 3655 14382
rect -3735 14222 -3655 14302
rect -3425 14222 -3345 14302
rect -1965 14222 -1885 14302
rect -1655 14222 -1575 14302
rect -195 14222 -115 14302
rect 115 14222 195 14302
rect 1575 14222 1655 14302
rect 1885 14222 1965 14302
rect 3345 14222 3425 14302
rect 3655 14222 3735 14302
rect -3735 11618 -3655 11698
rect -3425 11618 -3345 11698
rect -1965 11618 -1885 11698
rect -1655 11618 -1575 11698
rect -195 11618 -115 11698
rect 115 11618 195 11698
rect 1575 11618 1655 11698
rect 1885 11618 1965 11698
rect 3345 11618 3425 11698
rect 3655 11618 3735 11698
rect -3655 11538 -3575 11618
rect -3505 11538 -3425 11618
rect -1885 11538 -1805 11618
rect -1735 11538 -1655 11618
rect -115 11538 -35 11618
rect 35 11538 115 11618
rect 1655 11538 1735 11618
rect 1805 11538 1885 11618
rect 3425 11538 3505 11618
rect 3575 11538 3655 11618
rect -3005 10210 -2305 10280
rect -1235 10210 -535 10280
rect 535 10210 1235 10280
rect 2305 10210 3005 10280
rect -2770 10045 -2690 10125
rect -2620 10045 -2540 10125
rect -1000 10045 -920 10125
rect -850 10045 -770 10125
rect 770 10045 850 10125
rect 920 10045 1000 10125
rect 2540 10045 2620 10125
rect 2690 10045 2770 10125
rect -2850 9965 -2460 10045
rect -1080 9965 -690 10045
rect 690 9965 1080 10045
rect 2460 9965 2850 10045
rect -2825 9895 -2485 9965
rect -1055 9895 -715 9965
rect 715 9895 1055 9965
rect 2485 9895 2825 9965
rect -2850 9815 -2460 9895
rect -1080 9815 -690 9895
rect 690 9815 1080 9895
rect 2460 9815 2850 9895
rect -2770 9735 -2690 9815
rect -2620 9735 -2540 9815
rect -1000 9735 -920 9815
rect -850 9735 -770 9815
rect 770 9735 850 9815
rect 920 9735 1000 9815
rect 2540 9735 2620 9815
rect 2690 9735 2770 9815
rect -3655 7882 -3575 7962
rect -3505 7882 -3425 7962
rect -1885 7882 -1805 7962
rect -1735 7882 -1655 7962
rect -115 7882 -35 7962
rect 35 7882 115 7962
rect 1655 7882 1735 7962
rect 1805 7882 1885 7962
rect 3425 7882 3505 7962
rect 3575 7882 3655 7962
rect -3735 7802 -3655 7882
rect -3425 7802 -3345 7882
rect -1965 7802 -1885 7882
rect -1655 7802 -1575 7882
rect -195 7802 -115 7882
rect 115 7802 195 7882
rect 1575 7802 1655 7882
rect 1885 7802 1965 7882
rect 3345 7802 3425 7882
rect 3655 7802 3735 7882
rect -3735 5198 -3655 5278
rect -3425 5198 -3345 5278
rect -1965 5198 -1885 5278
rect -1655 5198 -1575 5278
rect -195 5198 -115 5278
rect 115 5198 195 5278
rect 1575 5198 1655 5278
rect 1885 5198 1965 5278
rect 3345 5198 3425 5278
rect 3655 5198 3735 5278
rect -3655 5118 -3575 5198
rect -3505 5118 -3425 5198
rect -1885 5118 -1805 5198
rect -1735 5118 -1655 5198
rect -115 5118 -35 5198
rect 35 5118 115 5198
rect 1655 5118 1735 5198
rect 1805 5118 1885 5198
rect 3425 5118 3505 5198
rect 3575 5118 3655 5198
rect -3005 3790 -2305 3860
rect -1235 3790 -535 3860
rect 535 3790 1235 3860
rect 2305 3790 3005 3860
rect -2770 3625 -2690 3705
rect -2620 3625 -2540 3705
rect -1000 3625 -920 3705
rect -850 3625 -770 3705
rect 770 3625 850 3705
rect 920 3625 1000 3705
rect 2540 3625 2620 3705
rect 2690 3625 2770 3705
rect -2850 3545 -2460 3625
rect -1080 3545 -690 3625
rect 690 3545 1080 3625
rect 2460 3545 2850 3625
rect -2825 3475 -2485 3545
rect -1055 3475 -715 3545
rect 715 3475 1055 3545
rect 2485 3475 2825 3545
rect -2850 3395 -2460 3475
rect -1080 3395 -690 3475
rect 690 3395 1080 3475
rect 2460 3395 2850 3475
rect -2770 3315 -2690 3395
rect -2620 3315 -2540 3395
rect -1000 3315 -920 3395
rect -850 3315 -770 3395
rect 770 3315 850 3395
rect 920 3315 1000 3395
rect 2540 3315 2620 3395
rect 2690 3315 2770 3395
rect -3655 1462 -3575 1542
rect -3505 1462 -3425 1542
rect -1885 1462 -1805 1542
rect -1735 1462 -1655 1542
rect -115 1462 -35 1542
rect 35 1462 115 1542
rect 1655 1462 1735 1542
rect 1805 1462 1885 1542
rect 3425 1462 3505 1542
rect 3575 1462 3655 1542
rect -3735 1382 -3655 1462
rect -3425 1382 -3345 1462
rect -1965 1382 -1885 1462
rect -1655 1382 -1575 1462
rect -195 1382 -115 1462
rect 115 1382 195 1462
rect 1575 1382 1655 1462
rect 1885 1382 1965 1462
rect 3345 1382 3425 1462
rect 3655 1382 3735 1462
rect -3735 -1222 -3655 -1142
rect -3425 -1222 -3345 -1142
rect -1965 -1222 -1885 -1142
rect -1655 -1222 -1575 -1142
rect -195 -1222 -115 -1142
rect 115 -1222 195 -1142
rect 1575 -1222 1655 -1142
rect 1885 -1222 1965 -1142
rect 3345 -1222 3425 -1142
rect 3655 -1222 3735 -1142
rect -3655 -1302 -3575 -1222
rect -3505 -1302 -3425 -1222
rect -1885 -1302 -1805 -1222
rect -1735 -1302 -1655 -1222
rect -115 -1302 -35 -1222
rect 35 -1302 115 -1222
rect 1655 -1302 1735 -1222
rect 1805 -1302 1885 -1222
rect 3425 -1302 3505 -1222
rect 3575 -1302 3655 -1222
rect -3005 -2630 -2305 -2560
rect -1235 -2630 -535 -2560
rect 535 -2630 1235 -2560
rect 2305 -2630 3005 -2560
rect -2770 -2795 -2690 -2715
rect -2620 -2795 -2540 -2715
rect -1000 -2795 -920 -2715
rect -850 -2795 -770 -2715
rect 770 -2795 850 -2715
rect 920 -2795 1000 -2715
rect 2540 -2795 2620 -2715
rect 2690 -2795 2770 -2715
rect -2850 -2875 -2460 -2795
rect -1080 -2875 -690 -2795
rect 690 -2875 1080 -2795
rect 2460 -2875 2850 -2795
rect -2825 -2945 -2485 -2875
rect -1055 -2945 -715 -2875
rect 715 -2945 1055 -2875
rect 2485 -2945 2825 -2875
rect -2850 -3025 -2460 -2945
rect -1080 -3025 -690 -2945
rect 690 -3025 1080 -2945
rect 2460 -3025 2850 -2945
rect -2770 -3105 -2690 -3025
rect -2620 -3105 -2540 -3025
rect -1000 -3105 -920 -3025
rect -850 -3105 -770 -3025
rect 770 -3105 850 -3025
rect 920 -3105 1000 -3025
rect 2540 -3105 2620 -3025
rect 2690 -3105 2770 -3025
rect -3655 -4958 -3575 -4878
rect -3505 -4958 -3425 -4878
rect -1885 -4958 -1805 -4878
rect -1735 -4958 -1655 -4878
rect -115 -4958 -35 -4878
rect 35 -4958 115 -4878
rect 1655 -4958 1735 -4878
rect 1805 -4958 1885 -4878
rect 3425 -4958 3505 -4878
rect 3575 -4958 3655 -4878
rect -3735 -5038 -3655 -4958
rect -3425 -5038 -3345 -4958
rect -1965 -5038 -1885 -4958
rect -1655 -5038 -1575 -4958
rect -195 -5038 -115 -4958
rect 115 -5038 195 -4958
rect 1575 -5038 1655 -4958
rect 1885 -5038 1965 -4958
rect 3345 -5038 3425 -4958
rect 3655 -5038 3735 -4958
rect -3735 -7642 -3655 -7562
rect -3425 -7642 -3345 -7562
rect -1965 -7642 -1885 -7562
rect -1655 -7642 -1575 -7562
rect -195 -7642 -115 -7562
rect 115 -7642 195 -7562
rect 1575 -7642 1655 -7562
rect 1885 -7642 1965 -7562
rect 3345 -7642 3425 -7562
rect 3655 -7642 3735 -7562
rect -3655 -7722 -3575 -7642
rect -3505 -7722 -3425 -7642
rect -1885 -7722 -1805 -7642
rect -1735 -7722 -1655 -7642
rect -115 -7722 -35 -7642
rect 35 -7722 115 -7642
rect 1655 -7722 1735 -7642
rect 1805 -7722 1885 -7642
rect 3425 -7722 3505 -7642
rect 3575 -7722 3655 -7642
rect -3005 -9050 -2305 -8980
rect -1235 -9050 -535 -8980
rect 535 -9050 1235 -8980
rect 2305 -9050 3005 -8980
rect -2770 -9215 -2690 -9135
rect -2620 -9215 -2540 -9135
rect -1000 -9215 -920 -9135
rect -850 -9215 -770 -9135
rect 770 -9215 850 -9135
rect 920 -9215 1000 -9135
rect 2540 -9215 2620 -9135
rect 2690 -9215 2770 -9135
rect -2850 -9295 -2460 -9215
rect -1080 -9295 -690 -9215
rect 690 -9295 1080 -9215
rect 2460 -9295 2850 -9215
rect -2825 -9365 -2485 -9295
rect -1055 -9365 -715 -9295
rect 715 -9365 1055 -9295
rect 2485 -9365 2825 -9295
rect -2850 -9445 -2460 -9365
rect -1080 -9445 -690 -9365
rect 690 -9445 1080 -9365
rect 2460 -9445 2850 -9365
rect -2770 -9525 -2690 -9445
rect -2620 -9525 -2540 -9445
rect -1000 -9525 -920 -9445
rect -850 -9525 -770 -9445
rect 770 -9525 850 -9445
rect 920 -9525 1000 -9445
rect 2540 -9525 2620 -9445
rect 2690 -9525 2770 -9445
rect -3655 -11378 -3575 -11298
rect -3505 -11378 -3425 -11298
rect -1885 -11378 -1805 -11298
rect -1735 -11378 -1655 -11298
rect -115 -11378 -35 -11298
rect 35 -11378 115 -11298
rect 1655 -11378 1735 -11298
rect 1805 -11378 1885 -11298
rect 3425 -11378 3505 -11298
rect 3575 -11378 3655 -11298
rect -3735 -11458 -3655 -11378
rect -3425 -11458 -3345 -11378
rect -1965 -11458 -1885 -11378
rect -1655 -11458 -1575 -11378
rect -195 -11458 -115 -11378
rect 115 -11458 195 -11378
rect 1575 -11458 1655 -11378
rect 1885 -11458 1965 -11378
rect 3345 -11458 3425 -11378
rect 3655 -11458 3735 -11378
rect -3735 -14062 -3655 -13982
rect -3425 -14062 -3345 -13982
rect -1965 -14062 -1885 -13982
rect -1655 -14062 -1575 -13982
rect -195 -14062 -115 -13982
rect 115 -14062 195 -13982
rect 1575 -14062 1655 -13982
rect 1885 -14062 1965 -13982
rect 3345 -14062 3425 -13982
rect 3655 -14062 3735 -13982
rect -3655 -14142 -3575 -14062
rect -3505 -14142 -3425 -14062
rect -1885 -14142 -1805 -14062
rect -1735 -14142 -1655 -14062
rect -115 -14142 -35 -14062
rect 35 -14142 115 -14062
rect 1655 -14142 1735 -14062
rect 1805 -14142 1885 -14062
rect 3425 -14142 3505 -14062
rect 3575 -14142 3655 -14062
rect -3005 -15470 -2305 -15400
rect -1235 -15470 -535 -15400
rect 535 -15470 1235 -15400
rect 2305 -15470 3005 -15400
rect -2770 -15635 -2690 -15555
rect -2620 -15635 -2540 -15555
rect -1000 -15635 -920 -15555
rect -850 -15635 -770 -15555
rect 770 -15635 850 -15555
rect 920 -15635 1000 -15555
rect 2540 -15635 2620 -15555
rect 2690 -15635 2770 -15555
rect -2850 -15715 -2460 -15635
rect -1080 -15715 -690 -15635
rect 690 -15715 1080 -15635
rect 2460 -15715 2850 -15635
rect -4425 -15820 -4345 -15740
rect -4115 -15820 -4035 -15740
rect -2825 -15785 -2485 -15715
rect -1055 -15785 -715 -15715
rect 715 -15785 1055 -15715
rect 2485 -15785 2825 -15715
rect 4350 -15740 4410 15740
rect -4410 -16340 -4350 -15820
rect -4345 -15900 -4265 -15820
rect -4195 -15900 -4115 -15820
rect -2850 -15865 -2460 -15785
rect -1080 -15865 -690 -15785
rect 690 -15865 1080 -15785
rect 2460 -15865 2850 -15785
rect 4035 -15820 4115 -15740
rect 4345 -15820 4425 -15740
rect -2770 -15945 -2690 -15865
rect -2620 -15945 -2540 -15865
rect -1000 -15945 -920 -15865
rect -850 -15945 -770 -15865
rect 770 -15945 850 -15865
rect 920 -15945 1000 -15865
rect 2540 -15945 2620 -15865
rect 2690 -15945 2770 -15865
rect 4115 -15900 4195 -15820
rect 4265 -15900 4345 -15820
rect 4350 -16340 4410 -15820
rect -4410 -16400 4410 -16340
rect 4530 -16520 4590 16520
rect -4590 -16580 4590 -16520
<< nwell >>
rect -4530 -16520 4530 16520
<< pmos >>
rect -3280 10210 -2030 15710
rect -1510 10210 -260 15710
rect 260 10210 1510 15710
rect 2030 10210 3280 15710
rect -3280 3790 -2030 9290
rect -1510 3790 -260 9290
rect 260 3790 1510 9290
rect 2030 3790 3280 9290
rect -3280 -2630 -2030 2870
rect -1510 -2630 -260 2870
rect 260 -2630 1510 2870
rect 2030 -2630 3280 2870
rect -3280 -9050 -2030 -3550
rect -1510 -9050 -260 -3550
rect 260 -9050 1510 -3550
rect 2030 -9050 3280 -3550
rect -3280 -15470 -2030 -9970
rect -1510 -15470 -260 -9970
rect 260 -15470 1510 -9970
rect 2030 -15470 3280 -9970
<< pdiff >>
rect -3655 14367 -3280 15710
rect -3720 14302 -3280 14367
rect -3720 11618 -3655 14302
rect -3425 11618 -3280 14302
rect -3720 11553 -3280 11618
rect -3655 10210 -3280 11553
rect -2030 14302 -1510 15710
rect -2030 11618 -1885 14302
rect -1655 11618 -1510 14302
rect -2030 10210 -1510 11618
rect -260 14302 260 15710
rect -260 11618 -115 14302
rect 115 11618 260 14302
rect -260 10210 260 11618
rect 1510 14302 2030 15710
rect 1510 11618 1655 14302
rect 1885 11618 2030 14302
rect 1510 10210 2030 11618
rect 3280 14367 3655 15710
rect 3280 14302 3720 14367
rect 3280 11618 3425 14302
rect 3655 11618 3720 14302
rect 3280 11553 3720 11618
rect 3280 10210 3655 11553
rect -3655 7947 -3280 9290
rect -3720 7882 -3280 7947
rect -3720 5198 -3655 7882
rect -3425 5198 -3280 7882
rect -3720 5133 -3280 5198
rect -3655 3790 -3280 5133
rect -2030 7882 -1510 9290
rect -2030 5198 -1885 7882
rect -1655 5198 -1510 7882
rect -2030 3790 -1510 5198
rect -260 7882 260 9290
rect -260 5198 -115 7882
rect 115 5198 260 7882
rect -260 3790 260 5198
rect 1510 7882 2030 9290
rect 1510 5198 1655 7882
rect 1885 5198 2030 7882
rect 1510 3790 2030 5198
rect 3280 7947 3655 9290
rect 3280 7882 3720 7947
rect 3280 5198 3425 7882
rect 3655 5198 3720 7882
rect 3280 5133 3720 5198
rect 3280 3790 3655 5133
rect -3655 1527 -3280 2870
rect -3720 1462 -3280 1527
rect -3720 -1222 -3655 1462
rect -3425 -1222 -3280 1462
rect -3720 -1287 -3280 -1222
rect -3655 -2630 -3280 -1287
rect -2030 1462 -1510 2870
rect -2030 -1222 -1885 1462
rect -1655 -1222 -1510 1462
rect -2030 -2630 -1510 -1222
rect -260 1462 260 2870
rect -260 -1222 -115 1462
rect 115 -1222 260 1462
rect -260 -2630 260 -1222
rect 1510 1462 2030 2870
rect 1510 -1222 1655 1462
rect 1885 -1222 2030 1462
rect 1510 -2630 2030 -1222
rect 3280 1527 3655 2870
rect 3280 1462 3720 1527
rect 3280 -1222 3425 1462
rect 3655 -1222 3720 1462
rect 3280 -1287 3720 -1222
rect 3280 -2630 3655 -1287
rect -3655 -4893 -3280 -3550
rect -3720 -4958 -3280 -4893
rect -3720 -7642 -3655 -4958
rect -3425 -7642 -3280 -4958
rect -3720 -7707 -3280 -7642
rect -3655 -9050 -3280 -7707
rect -2030 -4958 -1510 -3550
rect -2030 -7642 -1885 -4958
rect -1655 -7642 -1510 -4958
rect -2030 -9050 -1510 -7642
rect -260 -4958 260 -3550
rect -260 -7642 -115 -4958
rect 115 -7642 260 -4958
rect -260 -9050 260 -7642
rect 1510 -4958 2030 -3550
rect 1510 -7642 1655 -4958
rect 1885 -7642 2030 -4958
rect 1510 -9050 2030 -7642
rect 3280 -4893 3655 -3550
rect 3280 -4958 3720 -4893
rect 3280 -7642 3425 -4958
rect 3655 -7642 3720 -4958
rect 3280 -7707 3720 -7642
rect 3280 -9050 3655 -7707
rect -3655 -11313 -3280 -9970
rect -3720 -11378 -3280 -11313
rect -3720 -14062 -3655 -11378
rect -3425 -14062 -3280 -11378
rect -3720 -14127 -3280 -14062
rect -3655 -15470 -3280 -14127
rect -2030 -11378 -1510 -9970
rect -2030 -14062 -1885 -11378
rect -1655 -14062 -1510 -11378
rect -2030 -15470 -1510 -14062
rect -260 -11378 260 -9970
rect -260 -14062 -115 -11378
rect 115 -14062 260 -11378
rect -260 -15470 260 -14062
rect 1510 -11378 2030 -9970
rect 1510 -14062 1655 -11378
rect 1885 -14062 2030 -11378
rect 1510 -15470 2030 -14062
rect 3280 -11313 3655 -9970
rect 3280 -11378 3720 -11313
rect 3280 -14062 3425 -11378
rect 3655 -14062 3720 -11378
rect 3280 -14127 3720 -14062
rect 3280 -15470 3655 -14127
<< pdiffc >>
rect -3655 11618 -3425 14302
rect -1885 11618 -1655 14302
rect -115 11618 115 14302
rect 1655 11618 1885 14302
rect 3425 11618 3655 14302
rect -3655 5198 -3425 7882
rect -1885 5198 -1655 7882
rect -115 5198 115 7882
rect 1655 5198 1885 7882
rect 3425 5198 3655 7882
rect -3655 -1222 -3425 1462
rect -1885 -1222 -1655 1462
rect -115 -1222 115 1462
rect 1655 -1222 1885 1462
rect 3425 -1222 3655 1462
rect -3655 -7642 -3425 -4958
rect -1885 -7642 -1655 -4958
rect -115 -7642 115 -4958
rect 1655 -7642 1885 -4958
rect 3425 -7642 3655 -4958
rect -3655 -14062 -3425 -11378
rect -1885 -14062 -1655 -11378
rect -115 -14062 115 -11378
rect 1655 -14062 1885 -11378
rect 3425 -14062 3655 -11378
<< nsubdiff >>
rect -4410 16040 4410 16400
rect -4410 15820 -4050 16040
rect -4410 -15820 -4345 15820
rect -4115 -15820 -4050 15820
rect 4050 15820 4410 16040
rect -4410 -16040 -4050 -15820
rect 4050 -15820 4115 15820
rect 4345 -15820 4410 15820
rect 4050 -16040 4410 -15820
rect -4410 -16400 4410 -16040
<< nsubdiffcont >>
rect -4345 -15820 -4115 15820
rect 4115 -15820 4345 15820
<< poly >>
rect -3280 15710 -2030 15930
rect -1510 15710 -260 15930
rect 260 15710 1510 15930
rect 2030 15710 3280 15930
rect -3280 10045 -2030 10210
rect -3280 9930 -2770 10045
rect -2835 9815 -2770 9930
rect -2540 9930 -2030 10045
rect -1510 10045 -260 10210
rect -1510 9930 -1000 10045
rect -2540 9815 -2475 9930
rect -2835 9750 -2475 9815
rect -1065 9815 -1000 9930
rect -770 9930 -260 10045
rect 260 10045 1510 10210
rect 260 9930 770 10045
rect -770 9815 -705 9930
rect -1065 9750 -705 9815
rect 705 9815 770 9930
rect 1000 9930 1510 10045
rect 2030 10045 3280 10210
rect 2030 9930 2540 10045
rect 1000 9815 1065 9930
rect 705 9750 1065 9815
rect 2475 9815 2540 9930
rect 2770 9930 3280 10045
rect 2770 9815 2835 9930
rect 2475 9750 2835 9815
rect -3280 9290 -2030 9510
rect -1510 9290 -260 9510
rect 260 9290 1510 9510
rect 2030 9290 3280 9510
rect -3280 3625 -2030 3790
rect -3280 3510 -2770 3625
rect -2835 3395 -2770 3510
rect -2540 3510 -2030 3625
rect -1510 3625 -260 3790
rect -1510 3510 -1000 3625
rect -2540 3395 -2475 3510
rect -2835 3330 -2475 3395
rect -1065 3395 -1000 3510
rect -770 3510 -260 3625
rect 260 3625 1510 3790
rect 260 3510 770 3625
rect -770 3395 -705 3510
rect -1065 3330 -705 3395
rect 705 3395 770 3510
rect 1000 3510 1510 3625
rect 2030 3625 3280 3790
rect 2030 3510 2540 3625
rect 1000 3395 1065 3510
rect 705 3330 1065 3395
rect 2475 3395 2540 3510
rect 2770 3510 3280 3625
rect 2770 3395 2835 3510
rect 2475 3330 2835 3395
rect -3280 2870 -2030 3090
rect -1510 2870 -260 3090
rect 260 2870 1510 3090
rect 2030 2870 3280 3090
rect -3280 -2795 -2030 -2630
rect -3280 -2910 -2770 -2795
rect -2835 -3025 -2770 -2910
rect -2540 -2910 -2030 -2795
rect -1510 -2795 -260 -2630
rect -1510 -2910 -1000 -2795
rect -2540 -3025 -2475 -2910
rect -2835 -3090 -2475 -3025
rect -1065 -3025 -1000 -2910
rect -770 -2910 -260 -2795
rect 260 -2795 1510 -2630
rect 260 -2910 770 -2795
rect -770 -3025 -705 -2910
rect -1065 -3090 -705 -3025
rect 705 -3025 770 -2910
rect 1000 -2910 1510 -2795
rect 2030 -2795 3280 -2630
rect 2030 -2910 2540 -2795
rect 1000 -3025 1065 -2910
rect 705 -3090 1065 -3025
rect 2475 -3025 2540 -2910
rect 2770 -2910 3280 -2795
rect 2770 -3025 2835 -2910
rect 2475 -3090 2835 -3025
rect -3280 -3550 -2030 -3330
rect -1510 -3550 -260 -3330
rect 260 -3550 1510 -3330
rect 2030 -3550 3280 -3330
rect -3280 -9215 -2030 -9050
rect -3280 -9330 -2770 -9215
rect -2835 -9445 -2770 -9330
rect -2540 -9330 -2030 -9215
rect -1510 -9215 -260 -9050
rect -1510 -9330 -1000 -9215
rect -2540 -9445 -2475 -9330
rect -2835 -9510 -2475 -9445
rect -1065 -9445 -1000 -9330
rect -770 -9330 -260 -9215
rect 260 -9215 1510 -9050
rect 260 -9330 770 -9215
rect -770 -9445 -705 -9330
rect -1065 -9510 -705 -9445
rect 705 -9445 770 -9330
rect 1000 -9330 1510 -9215
rect 2030 -9215 3280 -9050
rect 2030 -9330 2540 -9215
rect 1000 -9445 1065 -9330
rect 705 -9510 1065 -9445
rect 2475 -9445 2540 -9330
rect 2770 -9330 3280 -9215
rect 2770 -9445 2835 -9330
rect 2475 -9510 2835 -9445
rect -3280 -9970 -2030 -9750
rect -1510 -9970 -260 -9750
rect 260 -9970 1510 -9750
rect 2030 -9970 3280 -9750
rect -3280 -15635 -2030 -15470
rect -3280 -15750 -2770 -15635
rect -2835 -15865 -2770 -15750
rect -2540 -15750 -2030 -15635
rect -1510 -15635 -260 -15470
rect -1510 -15750 -1000 -15635
rect -2540 -15865 -2475 -15750
rect -2835 -15930 -2475 -15865
rect -1065 -15865 -1000 -15750
rect -770 -15750 -260 -15635
rect 260 -15635 1510 -15470
rect 260 -15750 770 -15635
rect -770 -15865 -705 -15750
rect -1065 -15930 -705 -15865
rect 705 -15865 770 -15750
rect 1000 -15750 1510 -15635
rect 2030 -15635 3280 -15470
rect 2030 -15750 2540 -15635
rect 1000 -15865 1065 -15750
rect 705 -15930 1065 -15865
rect 2475 -15865 2540 -15750
rect 2770 -15750 3280 -15635
rect 2770 -15865 2835 -15750
rect 2475 -15930 2835 -15865
<< polycont >>
rect -2770 9815 -2540 10045
rect -1000 9815 -770 10045
rect 770 9815 1000 10045
rect 2540 9815 2770 10045
rect -2770 3395 -2540 3625
rect -1000 3395 -770 3625
rect 770 3395 1000 3625
rect 2540 3395 2770 3625
rect -2770 -3025 -2540 -2795
rect -1000 -3025 -770 -2795
rect 770 -3025 1000 -2795
rect 2540 -3025 2770 -2795
rect -2770 -9445 -2540 -9215
rect -1000 -9445 -770 -9215
rect 770 -9445 1000 -9215
rect 2540 -9445 2770 -9215
rect -2770 -15865 -2540 -15635
rect -1000 -15865 -770 -15635
rect 770 -15865 1000 -15635
rect 2540 -15865 2770 -15635
<< metal1 >>
rect -4345 16105 4345 16335
rect -4345 -16105 -4115 16105
rect -3655 11563 -3425 14357
rect -1885 11563 -1655 14357
rect -115 11563 115 14357
rect 1655 11563 1885 14357
rect 3425 11563 3655 14357
rect -2825 9815 -2485 10045
rect -1055 9815 -715 10045
rect 715 9815 1055 10045
rect 2485 9815 2825 10045
rect -3655 5143 -3425 7937
rect -1885 5143 -1655 7937
rect -115 5143 115 7937
rect 1655 5143 1885 7937
rect 3425 5143 3655 7937
rect -2825 3395 -2485 3625
rect -1055 3395 -715 3625
rect 715 3395 1055 3625
rect 2485 3395 2825 3625
rect -3655 -1277 -3425 1517
rect -1885 -1277 -1655 1517
rect -115 -1277 115 1517
rect 1655 -1277 1885 1517
rect 3425 -1277 3655 1517
rect -2825 -3025 -2485 -2795
rect -1055 -3025 -715 -2795
rect 715 -3025 1055 -2795
rect 2485 -3025 2825 -2795
rect -3655 -7697 -3425 -4903
rect -1885 -7697 -1655 -4903
rect -115 -7697 115 -4903
rect 1655 -7697 1885 -4903
rect 3425 -7697 3655 -4903
rect -2825 -9445 -2485 -9215
rect -1055 -9445 -715 -9215
rect 715 -9445 1055 -9215
rect 2485 -9445 2825 -9215
rect -3655 -14117 -3425 -11323
rect -1885 -14117 -1655 -11323
rect -115 -14117 115 -11323
rect 1655 -14117 1885 -11323
rect 3425 -14117 3655 -11323
rect -2825 -15865 -2485 -15635
rect -1055 -15865 -715 -15635
rect 715 -15865 1055 -15635
rect 2485 -15865 2825 -15635
rect 4115 -16105 4345 16105
rect -4345 -16335 4345 -16105
<< properties >>
string FIXED_BBOX -4230 -16220 4230 16220
string gencell pfet_03v3
string library gf180mcu
string parameters w 5.5 l 1.25 m 5 nf 4 diffcov 50 polycov 20 guard 1 glc 1 grc 1 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 class mosfet full_metal 1 compatible {pfet_03v3 pfet_06v0}
<< end >>

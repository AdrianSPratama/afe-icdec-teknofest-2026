magic
tech sky130A
magscale 1 2
timestamp 1771116256
<< nwell >>
rect -1399 -528 1399 528
<< pmos >>
rect -1203 -380 -953 308
rect -895 -380 -645 308
rect -587 -380 -337 308
rect -279 -380 -29 308
rect 29 -380 279 308
rect 337 -380 587 308
rect 645 -380 895 308
rect 953 -380 1203 308
<< pdiff >>
rect -1261 296 -1203 308
rect -1261 -368 -1249 296
rect -1215 -368 -1203 296
rect -1261 -380 -1203 -368
rect -953 296 -895 308
rect -953 -368 -941 296
rect -907 -368 -895 296
rect -953 -380 -895 -368
rect -645 296 -587 308
rect -645 -368 -633 296
rect -599 -368 -587 296
rect -645 -380 -587 -368
rect -337 296 -279 308
rect -337 -368 -325 296
rect -291 -368 -279 296
rect -337 -380 -279 -368
rect -29 296 29 308
rect -29 -368 -17 296
rect 17 -368 29 296
rect -29 -380 29 -368
rect 279 296 337 308
rect 279 -368 291 296
rect 325 -368 337 296
rect 279 -380 337 -368
rect 587 296 645 308
rect 587 -368 599 296
rect 633 -368 645 296
rect 587 -380 645 -368
rect 895 296 953 308
rect 895 -368 907 296
rect 941 -368 953 296
rect 895 -380 953 -368
rect 1203 296 1261 308
rect 1203 -368 1215 296
rect 1249 -368 1261 296
rect 1203 -380 1261 -368
<< pdiffc >>
rect -1249 -368 -1215 296
rect -941 -368 -907 296
rect -633 -368 -599 296
rect -325 -368 -291 296
rect -17 -368 17 296
rect 291 -368 325 296
rect 599 -368 633 296
rect 907 -368 941 296
rect 1215 -368 1249 296
<< nsubdiff >>
rect -1363 458 -1267 492
rect 1267 458 1363 492
rect -1363 395 -1329 458
rect 1329 395 1363 458
rect -1363 -458 -1329 -395
rect 1329 -458 1363 -395
rect -1363 -492 -1267 -458
rect 1267 -492 1363 -458
<< nsubdiffcont >>
rect -1267 458 1267 492
rect -1363 -395 -1329 395
rect 1329 -395 1363 395
rect -1267 -492 1267 -458
<< poly >>
rect -1203 389 -953 405
rect -1203 355 -1187 389
rect -969 355 -953 389
rect -1203 308 -953 355
rect -895 389 -645 405
rect -895 355 -879 389
rect -661 355 -645 389
rect -895 308 -645 355
rect -587 389 -337 405
rect -587 355 -571 389
rect -353 355 -337 389
rect -587 308 -337 355
rect -279 389 -29 405
rect -279 355 -263 389
rect -45 355 -29 389
rect -279 308 -29 355
rect 29 389 279 405
rect 29 355 45 389
rect 263 355 279 389
rect 29 308 279 355
rect 337 389 587 405
rect 337 355 353 389
rect 571 355 587 389
rect 337 308 587 355
rect 645 389 895 405
rect 645 355 661 389
rect 879 355 895 389
rect 645 308 895 355
rect 953 389 1203 405
rect 953 355 969 389
rect 1187 355 1203 389
rect 953 308 1203 355
rect -1203 -406 -953 -380
rect -895 -406 -645 -380
rect -587 -406 -337 -380
rect -279 -406 -29 -380
rect 29 -406 279 -380
rect 337 -406 587 -380
rect 645 -406 895 -380
rect 953 -406 1203 -380
<< polycont >>
rect -1187 355 -969 389
rect -879 355 -661 389
rect -571 355 -353 389
rect -263 355 -45 389
rect 45 355 263 389
rect 353 355 571 389
rect 661 355 879 389
rect 969 355 1187 389
<< locali >>
rect -1363 458 -1267 492
rect 1267 458 1363 492
rect -1363 395 -1329 458
rect 1329 395 1363 458
rect -1203 355 -1187 389
rect -969 355 -953 389
rect -895 355 -879 389
rect -661 355 -645 389
rect -587 355 -571 389
rect -353 355 -337 389
rect -279 355 -263 389
rect -45 355 -29 389
rect 29 355 45 389
rect 263 355 279 389
rect 337 355 353 389
rect 571 355 587 389
rect 645 355 661 389
rect 879 355 895 389
rect 953 355 969 389
rect 1187 355 1203 389
rect -1249 296 -1215 312
rect -1249 -384 -1215 -368
rect -941 296 -907 312
rect -941 -384 -907 -368
rect -633 296 -599 312
rect -633 -384 -599 -368
rect -325 296 -291 312
rect -325 -384 -291 -368
rect -17 296 17 312
rect -17 -384 17 -368
rect 291 296 325 312
rect 291 -384 325 -368
rect 599 296 633 312
rect 599 -384 633 -368
rect 907 296 941 312
rect 907 -384 941 -368
rect 1215 296 1249 312
rect 1215 -384 1249 -368
rect -1363 -458 -1329 -395
rect 1329 -458 1363 -395
rect -1363 -492 -1267 -458
rect 1267 -492 1363 -458
<< viali >>
rect -1187 355 -969 389
rect -879 355 -661 389
rect -571 355 -353 389
rect -263 355 -45 389
rect 45 355 263 389
rect 353 355 571 389
rect 661 355 879 389
rect 969 355 1187 389
rect -1249 -368 -1215 296
rect -941 -368 -907 296
rect -633 -368 -599 296
rect -325 -368 -291 296
rect -17 -368 17 296
rect 291 -368 325 296
rect 599 -368 633 296
rect 907 -368 941 296
rect 1215 -368 1249 296
<< metal1 >>
rect -1199 389 -957 395
rect -1199 355 -1187 389
rect -969 355 -957 389
rect -1199 349 -957 355
rect -891 389 -649 395
rect -891 355 -879 389
rect -661 355 -649 389
rect -891 349 -649 355
rect -583 389 -341 395
rect -583 355 -571 389
rect -353 355 -341 389
rect -583 349 -341 355
rect -275 389 -33 395
rect -275 355 -263 389
rect -45 355 -33 389
rect -275 349 -33 355
rect 33 389 275 395
rect 33 355 45 389
rect 263 355 275 389
rect 33 349 275 355
rect 341 389 583 395
rect 341 355 353 389
rect 571 355 583 389
rect 341 349 583 355
rect 649 389 891 395
rect 649 355 661 389
rect 879 355 891 389
rect 649 349 891 355
rect 957 389 1199 395
rect 957 355 969 389
rect 1187 355 1199 389
rect 957 349 1199 355
rect -1255 296 -1209 308
rect -1255 -368 -1249 296
rect -1215 -368 -1209 296
rect -1255 -380 -1209 -368
rect -947 296 -901 308
rect -947 -368 -941 296
rect -907 -368 -901 296
rect -947 -380 -901 -368
rect -639 296 -593 308
rect -639 -368 -633 296
rect -599 -368 -593 296
rect -639 -380 -593 -368
rect -331 296 -285 308
rect -331 -368 -325 296
rect -291 -368 -285 296
rect -331 -380 -285 -368
rect -23 296 23 308
rect -23 -368 -17 296
rect 17 -368 23 296
rect -23 -380 23 -368
rect 285 296 331 308
rect 285 -368 291 296
rect 325 -368 331 296
rect 285 -380 331 -368
rect 593 296 639 308
rect 593 -368 599 296
rect 633 -368 639 296
rect 593 -380 639 -368
rect 901 296 947 308
rect 901 -368 907 296
rect 941 -368 947 296
rect 901 -380 947 -368
rect 1209 296 1255 308
rect 1209 -368 1215 296
rect 1249 -368 1255 296
rect 1209 -380 1255 -368
<< properties >>
string FIXED_BBOX -1346 -475 1346 475
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 3.4375 l 1.25 m 1 nf 8 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 class mosfet compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1770979109
<< nwell >>
rect -2283 -719 2283 719
<< pmos >>
rect -2087 -500 -1087 500
rect -1029 -500 -29 500
rect 29 -500 1029 500
rect 1087 -500 2087 500
<< pdiff >>
rect -2145 488 -2087 500
rect -2145 -488 -2133 488
rect -2099 -488 -2087 488
rect -2145 -500 -2087 -488
rect -1087 488 -1029 500
rect -1087 -488 -1075 488
rect -1041 -488 -1029 488
rect -1087 -500 -1029 -488
rect -29 488 29 500
rect -29 -488 -17 488
rect 17 -488 29 488
rect -29 -500 29 -488
rect 1029 488 1087 500
rect 1029 -488 1041 488
rect 1075 -488 1087 488
rect 1029 -500 1087 -488
rect 2087 488 2145 500
rect 2087 -488 2099 488
rect 2133 -488 2145 488
rect 2087 -500 2145 -488
<< pdiffc >>
rect -2133 -488 -2099 488
rect -1075 -488 -1041 488
rect -17 -488 17 488
rect 1041 -488 1075 488
rect 2099 -488 2133 488
<< nsubdiff >>
rect -2247 649 -2151 683
rect 2151 649 2247 683
rect -2247 587 -2213 649
rect 2213 587 2247 649
rect -2247 -649 -2213 -587
rect 2213 -649 2247 -587
rect -2247 -683 -2151 -649
rect 2151 -683 2247 -649
<< nsubdiffcont >>
rect -2151 649 2151 683
rect -2247 -587 -2213 587
rect 2213 -587 2247 587
rect -2151 -683 2151 -649
<< poly >>
rect -2087 581 -1087 597
rect -2087 547 -2071 581
rect -1103 547 -1087 581
rect -2087 500 -1087 547
rect -1029 581 -29 597
rect -1029 547 -1013 581
rect -45 547 -29 581
rect -1029 500 -29 547
rect 29 581 1029 597
rect 29 547 45 581
rect 1013 547 1029 581
rect 29 500 1029 547
rect 1087 581 2087 597
rect 1087 547 1103 581
rect 2071 547 2087 581
rect 1087 500 2087 547
rect -2087 -547 -1087 -500
rect -2087 -581 -2071 -547
rect -1103 -581 -1087 -547
rect -2087 -597 -1087 -581
rect -1029 -547 -29 -500
rect -1029 -581 -1013 -547
rect -45 -581 -29 -547
rect -1029 -597 -29 -581
rect 29 -547 1029 -500
rect 29 -581 45 -547
rect 1013 -581 1029 -547
rect 29 -597 1029 -581
rect 1087 -547 2087 -500
rect 1087 -581 1103 -547
rect 2071 -581 2087 -547
rect 1087 -597 2087 -581
<< polycont >>
rect -2071 547 -1103 581
rect -1013 547 -45 581
rect 45 547 1013 581
rect 1103 547 2071 581
rect -2071 -581 -1103 -547
rect -1013 -581 -45 -547
rect 45 -581 1013 -547
rect 1103 -581 2071 -547
<< locali >>
rect -2247 649 -2151 683
rect 2151 649 2247 683
rect -2247 587 -2213 649
rect 2213 587 2247 649
rect -2087 547 -2071 581
rect -1103 547 -1087 581
rect -1029 547 -1013 581
rect -45 547 -29 581
rect 29 547 45 581
rect 1013 547 1029 581
rect 1087 547 1103 581
rect 2071 547 2087 581
rect -2133 488 -2099 504
rect -2133 -504 -2099 -488
rect -1075 488 -1041 504
rect -1075 -504 -1041 -488
rect -17 488 17 504
rect -17 -504 17 -488
rect 1041 488 1075 504
rect 1041 -504 1075 -488
rect 2099 488 2133 504
rect 2099 -504 2133 -488
rect -2087 -581 -2071 -547
rect -1103 -581 -1087 -547
rect -1029 -581 -1013 -547
rect -45 -581 -29 -547
rect 29 -581 45 -547
rect 1013 -581 1029 -547
rect 1087 -581 1103 -547
rect 2071 -581 2087 -547
rect -2247 -649 -2213 -587
rect 2213 -649 2247 -587
rect -2247 -683 -2151 -649
rect 2151 -683 2247 -649
<< viali >>
rect -2071 547 -1103 581
rect -1013 547 -45 581
rect 45 547 1013 581
rect 1103 547 2071 581
rect -2133 -488 -2099 488
rect -1075 -488 -1041 488
rect -17 -488 17 488
rect 1041 -488 1075 488
rect 2099 -488 2133 488
rect -2071 -581 -1103 -547
rect -1013 -581 -45 -547
rect 45 -581 1013 -547
rect 1103 -581 2071 -547
<< metal1 >>
rect -2083 581 -1091 587
rect -2083 547 -2071 581
rect -1103 547 -1091 581
rect -2083 541 -1091 547
rect -1025 581 -33 587
rect -1025 547 -1013 581
rect -45 547 -33 581
rect -1025 541 -33 547
rect 33 581 1025 587
rect 33 547 45 581
rect 1013 547 1025 581
rect 33 541 1025 547
rect 1091 581 2083 587
rect 1091 547 1103 581
rect 2071 547 2083 581
rect 1091 541 2083 547
rect -2139 488 -2093 500
rect -2139 -488 -2133 488
rect -2099 -488 -2093 488
rect -2139 -500 -2093 -488
rect -1081 488 -1035 500
rect -1081 -488 -1075 488
rect -1041 -488 -1035 488
rect -1081 -500 -1035 -488
rect -23 488 23 500
rect -23 -488 -17 488
rect 17 -488 23 488
rect -23 -500 23 -488
rect 1035 488 1081 500
rect 1035 -488 1041 488
rect 1075 -488 1081 488
rect 1035 -500 1081 -488
rect 2093 488 2139 500
rect 2093 -488 2099 488
rect 2133 -488 2139 488
rect 2093 -500 2139 -488
rect -2083 -547 -1091 -541
rect -2083 -581 -2071 -547
rect -1103 -581 -1091 -547
rect -2083 -587 -1091 -581
rect -1025 -547 -33 -541
rect -1025 -581 -1013 -547
rect -45 -581 -33 -547
rect -1025 -587 -33 -581
rect 33 -547 1025 -541
rect 33 -581 45 -547
rect 1013 -581 1025 -547
rect 33 -587 1025 -581
rect 1091 -547 2083 -541
rect 1091 -581 1103 -547
rect 2071 -581 2083 -547
rect 1091 -587 2083 -581
<< properties >>
string FIXED_BBOX -2230 -666 2230 666
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 5.0 l 5.0 m 1 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 class mosfet compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0 ad {int((nf+1)/2) * W/nf * 0.29} as {int((nf+2)/2) * W/nf * 0.29} pd {2*int((nf+1)/2) * (W/nf + 0.29)} ps {2*int((nf+2)/2) * (W/nf + 0.29)} nrd {0.29 / W} nrs {0.29 / W} sa 0 sb 0 sd 0 mult 1
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1771462974
<< error_p >>
rect -491 3125 -433 3131
rect -183 3125 -125 3131
rect 125 3125 183 3131
rect 433 3125 491 3131
rect -491 3091 -479 3125
rect -183 3091 -171 3125
rect 125 3091 137 3125
rect 433 3091 445 3125
rect -491 3085 -433 3091
rect -183 3085 -125 3091
rect 125 3085 183 3091
rect 433 3085 491 3091
rect -681 1882 681 2133
rect -491 1860 -433 1866
rect -183 1860 -125 1866
rect 125 1860 183 1866
rect 433 1860 491 1866
rect -491 1826 -479 1860
rect -183 1826 -171 1860
rect 125 1826 137 1860
rect 433 1826 445 1860
rect -491 1820 -433 1826
rect -183 1820 -125 1826
rect 125 1820 183 1826
rect 433 1820 491 1826
rect -681 617 681 868
rect -491 595 -433 601
rect -183 595 -125 601
rect 125 595 183 601
rect 433 595 491 601
rect -491 561 -479 595
rect -183 561 -171 595
rect 125 561 137 595
rect 433 561 445 595
rect -491 555 -433 561
rect -183 555 -125 561
rect 125 555 183 561
rect 433 555 491 561
rect -681 -648 681 -397
rect -491 -670 -433 -664
rect -183 -670 -125 -664
rect 125 -670 183 -664
rect 433 -670 491 -664
rect -491 -704 -479 -670
rect -183 -704 -171 -670
rect 125 -704 137 -670
rect 433 -704 445 -670
rect -491 -710 -433 -704
rect -183 -710 -125 -704
rect 125 -710 183 -704
rect 433 -710 491 -704
rect -681 -1913 681 -1662
rect -491 -1935 -433 -1929
rect -183 -1935 -125 -1929
rect 125 -1935 183 -1929
rect 433 -1935 491 -1929
rect -491 -1969 -479 -1935
rect -183 -1969 -171 -1935
rect 125 -1969 137 -1935
rect 433 -1969 445 -1935
rect -491 -1975 -433 -1969
rect -183 -1975 -125 -1969
rect 125 -1975 183 -1969
rect 433 -1975 491 -1969
<< nwell >>
rect -681 1882 681 3144
rect -681 617 681 1879
rect -681 -648 681 614
rect -681 -1913 681 -651
rect -681 -3178 681 -1916
<< pmos >>
rect -587 1944 -337 3044
rect -279 1944 -29 3044
rect 29 1944 279 3044
rect 337 1944 587 3044
rect -587 679 -337 1779
rect -279 679 -29 1779
rect 29 679 279 1779
rect 337 679 587 1779
rect -587 -586 -337 514
rect -279 -586 -29 514
rect 29 -586 279 514
rect 337 -586 587 514
rect -587 -1851 -337 -751
rect -279 -1851 -29 -751
rect 29 -1851 279 -751
rect 337 -1851 587 -751
rect -587 -3116 -337 -2016
rect -279 -3116 -29 -2016
rect 29 -3116 279 -2016
rect 337 -3116 587 -2016
<< pdiff >>
rect -645 2763 -587 3044
rect -645 2225 -633 2763
rect -599 2225 -587 2763
rect -645 1944 -587 2225
rect -337 2763 -279 3044
rect -337 2225 -325 2763
rect -291 2225 -279 2763
rect -337 1944 -279 2225
rect -29 2763 29 3044
rect -29 2225 -17 2763
rect 17 2225 29 2763
rect -29 1944 29 2225
rect 279 2763 337 3044
rect 279 2225 291 2763
rect 325 2225 337 2763
rect 279 1944 337 2225
rect 587 2763 645 3044
rect 587 2225 599 2763
rect 633 2225 645 2763
rect 587 1944 645 2225
rect -645 1498 -587 1779
rect -645 960 -633 1498
rect -599 960 -587 1498
rect -645 679 -587 960
rect -337 1498 -279 1779
rect -337 960 -325 1498
rect -291 960 -279 1498
rect -337 679 -279 960
rect -29 1498 29 1779
rect -29 960 -17 1498
rect 17 960 29 1498
rect -29 679 29 960
rect 279 1498 337 1779
rect 279 960 291 1498
rect 325 960 337 1498
rect 279 679 337 960
rect 587 1498 645 1779
rect 587 960 599 1498
rect 633 960 645 1498
rect 587 679 645 960
rect -645 233 -587 514
rect -645 -305 -633 233
rect -599 -305 -587 233
rect -645 -586 -587 -305
rect -337 233 -279 514
rect -337 -305 -325 233
rect -291 -305 -279 233
rect -337 -586 -279 -305
rect -29 233 29 514
rect -29 -305 -17 233
rect 17 -305 29 233
rect -29 -586 29 -305
rect 279 233 337 514
rect 279 -305 291 233
rect 325 -305 337 233
rect 279 -586 337 -305
rect 587 233 645 514
rect 587 -305 599 233
rect 633 -305 645 233
rect 587 -586 645 -305
rect -645 -1032 -587 -751
rect -645 -1570 -633 -1032
rect -599 -1570 -587 -1032
rect -645 -1851 -587 -1570
rect -337 -1032 -279 -751
rect -337 -1570 -325 -1032
rect -291 -1570 -279 -1032
rect -337 -1851 -279 -1570
rect -29 -1032 29 -751
rect -29 -1570 -17 -1032
rect 17 -1570 29 -1032
rect -29 -1851 29 -1570
rect 279 -1032 337 -751
rect 279 -1570 291 -1032
rect 325 -1570 337 -1032
rect 279 -1851 337 -1570
rect 587 -1032 645 -751
rect 587 -1570 599 -1032
rect 633 -1570 645 -1032
rect 587 -1851 645 -1570
rect -645 -2297 -587 -2016
rect -645 -2835 -633 -2297
rect -599 -2835 -587 -2297
rect -645 -3116 -587 -2835
rect -337 -2297 -279 -2016
rect -337 -2835 -325 -2297
rect -291 -2835 -279 -2297
rect -337 -3116 -279 -2835
rect -29 -2297 29 -2016
rect -29 -2835 -17 -2297
rect 17 -2835 29 -2297
rect -29 -3116 29 -2835
rect 279 -2297 337 -2016
rect 279 -2835 291 -2297
rect 325 -2835 337 -2297
rect 279 -3116 337 -2835
rect 587 -2297 645 -2016
rect 587 -2835 599 -2297
rect 633 -2835 645 -2297
rect 587 -3116 645 -2835
<< pdiffc >>
rect -633 2225 -599 2763
rect -325 2225 -291 2763
rect -17 2225 17 2763
rect 291 2225 325 2763
rect 599 2225 633 2763
rect -633 960 -599 1498
rect -325 960 -291 1498
rect -17 960 17 1498
rect 291 960 325 1498
rect 599 960 633 1498
rect -633 -305 -599 233
rect -325 -305 -291 233
rect -17 -305 17 233
rect 291 -305 325 233
rect 599 -305 633 233
rect -633 -1570 -599 -1032
rect -325 -1570 -291 -1032
rect -17 -1570 17 -1032
rect 291 -1570 325 -1032
rect 599 -1570 633 -1032
rect -633 -2835 -599 -2297
rect -325 -2835 -291 -2297
rect -17 -2835 17 -2297
rect 291 -2835 325 -2297
rect 599 -2835 633 -2297
<< poly >>
rect -500 3125 -424 3141
rect -500 3108 -484 3125
rect -587 3091 -484 3108
rect -440 3108 -424 3125
rect -192 3125 -116 3141
rect -192 3108 -176 3125
rect -440 3091 -337 3108
rect -587 3044 -337 3091
rect -279 3091 -176 3108
rect -132 3108 -116 3125
rect 116 3125 192 3141
rect 116 3108 132 3125
rect -132 3091 -29 3108
rect -279 3044 -29 3091
rect 29 3091 132 3108
rect 176 3108 192 3125
rect 424 3125 500 3141
rect 424 3108 440 3125
rect 176 3091 279 3108
rect 29 3044 279 3091
rect 337 3091 440 3108
rect 484 3108 500 3125
rect 484 3091 587 3108
rect 337 3044 587 3091
rect -587 1918 -337 1944
rect -279 1918 -29 1944
rect 29 1918 279 1944
rect 337 1918 587 1944
rect -500 1860 -424 1876
rect -500 1843 -484 1860
rect -587 1826 -484 1843
rect -440 1843 -424 1860
rect -192 1860 -116 1876
rect -192 1843 -176 1860
rect -440 1826 -337 1843
rect -587 1779 -337 1826
rect -279 1826 -176 1843
rect -132 1843 -116 1860
rect 116 1860 192 1876
rect 116 1843 132 1860
rect -132 1826 -29 1843
rect -279 1779 -29 1826
rect 29 1826 132 1843
rect 176 1843 192 1860
rect 424 1860 500 1876
rect 424 1843 440 1860
rect 176 1826 279 1843
rect 29 1779 279 1826
rect 337 1826 440 1843
rect 484 1843 500 1860
rect 484 1826 587 1843
rect 337 1779 587 1826
rect -587 653 -337 679
rect -279 653 -29 679
rect 29 653 279 679
rect 337 653 587 679
rect -500 595 -424 611
rect -500 578 -484 595
rect -587 561 -484 578
rect -440 578 -424 595
rect -192 595 -116 611
rect -192 578 -176 595
rect -440 561 -337 578
rect -587 514 -337 561
rect -279 561 -176 578
rect -132 578 -116 595
rect 116 595 192 611
rect 116 578 132 595
rect -132 561 -29 578
rect -279 514 -29 561
rect 29 561 132 578
rect 176 578 192 595
rect 424 595 500 611
rect 424 578 440 595
rect 176 561 279 578
rect 29 514 279 561
rect 337 561 440 578
rect 484 578 500 595
rect 484 561 587 578
rect 337 514 587 561
rect -587 -612 -337 -586
rect -279 -612 -29 -586
rect 29 -612 279 -586
rect 337 -612 587 -586
rect -500 -670 -424 -654
rect -500 -687 -484 -670
rect -587 -704 -484 -687
rect -440 -687 -424 -670
rect -192 -670 -116 -654
rect -192 -687 -176 -670
rect -440 -704 -337 -687
rect -587 -751 -337 -704
rect -279 -704 -176 -687
rect -132 -687 -116 -670
rect 116 -670 192 -654
rect 116 -687 132 -670
rect -132 -704 -29 -687
rect -279 -751 -29 -704
rect 29 -704 132 -687
rect 176 -687 192 -670
rect 424 -670 500 -654
rect 424 -687 440 -670
rect 176 -704 279 -687
rect 29 -751 279 -704
rect 337 -704 440 -687
rect 484 -687 500 -670
rect 484 -704 587 -687
rect 337 -751 587 -704
rect -587 -1877 -337 -1851
rect -279 -1877 -29 -1851
rect 29 -1877 279 -1851
rect 337 -1877 587 -1851
rect -500 -1935 -424 -1919
rect -500 -1952 -484 -1935
rect -587 -1969 -484 -1952
rect -440 -1952 -424 -1935
rect -192 -1935 -116 -1919
rect -192 -1952 -176 -1935
rect -440 -1969 -337 -1952
rect -587 -2016 -337 -1969
rect -279 -1969 -176 -1952
rect -132 -1952 -116 -1935
rect 116 -1935 192 -1919
rect 116 -1952 132 -1935
rect -132 -1969 -29 -1952
rect -279 -2016 -29 -1969
rect 29 -1969 132 -1952
rect 176 -1952 192 -1935
rect 424 -1935 500 -1919
rect 424 -1952 440 -1935
rect 176 -1969 279 -1952
rect 29 -2016 279 -1969
rect 337 -1969 440 -1952
rect 484 -1952 500 -1935
rect 484 -1969 587 -1952
rect 337 -2016 587 -1969
rect -587 -3142 -337 -3116
rect -279 -3142 -29 -3116
rect 29 -3142 279 -3116
rect 337 -3142 587 -3116
<< polycont >>
rect -484 3091 -440 3125
rect -176 3091 -132 3125
rect 132 3091 176 3125
rect 440 3091 484 3125
rect -484 1826 -440 1860
rect -176 1826 -132 1860
rect 132 1826 176 1860
rect 440 1826 484 1860
rect -484 561 -440 595
rect -176 561 -132 595
rect 132 561 176 595
rect 440 561 484 595
rect -484 -704 -440 -670
rect -176 -704 -132 -670
rect 132 -704 176 -670
rect 440 -704 484 -670
rect -484 -1969 -440 -1935
rect -176 -1969 -132 -1935
rect 132 -1969 176 -1935
rect 440 -1969 484 -1935
<< locali >>
rect -500 3091 -484 3125
rect -440 3091 -424 3125
rect -192 3091 -176 3125
rect -132 3091 -116 3125
rect 116 3091 132 3125
rect 176 3091 192 3125
rect 424 3091 440 3125
rect 484 3091 500 3125
rect -633 2763 -599 2779
rect -633 2209 -599 2225
rect -325 2763 -291 2779
rect -325 2209 -291 2225
rect -17 2763 17 2779
rect -17 2209 17 2225
rect 291 2763 325 2779
rect 291 2209 325 2225
rect 599 2763 633 2779
rect 599 2209 633 2225
rect -500 1826 -484 1860
rect -440 1826 -424 1860
rect -192 1826 -176 1860
rect -132 1826 -116 1860
rect 116 1826 132 1860
rect 176 1826 192 1860
rect 424 1826 440 1860
rect 484 1826 500 1860
rect -633 1498 -599 1514
rect -633 944 -599 960
rect -325 1498 -291 1514
rect -325 944 -291 960
rect -17 1498 17 1514
rect -17 944 17 960
rect 291 1498 325 1514
rect 291 944 325 960
rect 599 1498 633 1514
rect 599 944 633 960
rect -500 561 -484 595
rect -440 561 -424 595
rect -192 561 -176 595
rect -132 561 -116 595
rect 116 561 132 595
rect 176 561 192 595
rect 424 561 440 595
rect 484 561 500 595
rect -633 233 -599 249
rect -633 -321 -599 -305
rect -325 233 -291 249
rect -325 -321 -291 -305
rect -17 233 17 249
rect -17 -321 17 -305
rect 291 233 325 249
rect 291 -321 325 -305
rect 599 233 633 249
rect 599 -321 633 -305
rect -500 -704 -484 -670
rect -440 -704 -424 -670
rect -192 -704 -176 -670
rect -132 -704 -116 -670
rect 116 -704 132 -670
rect 176 -704 192 -670
rect 424 -704 440 -670
rect 484 -704 500 -670
rect -633 -1032 -599 -1016
rect -633 -1586 -599 -1570
rect -325 -1032 -291 -1016
rect -325 -1586 -291 -1570
rect -17 -1032 17 -1016
rect -17 -1586 17 -1570
rect 291 -1032 325 -1016
rect 291 -1586 325 -1570
rect 599 -1032 633 -1016
rect 599 -1586 633 -1570
rect -500 -1969 -484 -1935
rect -440 -1969 -424 -1935
rect -192 -1969 -176 -1935
rect -132 -1969 -116 -1935
rect 116 -1969 132 -1935
rect 176 -1969 192 -1935
rect 424 -1969 440 -1935
rect 484 -1969 500 -1935
rect -633 -2297 -599 -2281
rect -633 -2851 -599 -2835
rect -325 -2297 -291 -2281
rect -325 -2851 -291 -2835
rect -17 -2297 17 -2281
rect -17 -2851 17 -2835
rect 291 -2297 325 -2281
rect 291 -2851 325 -2835
rect 599 -2297 633 -2281
rect 599 -2851 633 -2835
<< viali >>
rect -479 3091 -445 3125
rect -171 3091 -137 3125
rect 137 3091 171 3125
rect 445 3091 479 3125
rect -633 2225 -599 2763
rect -325 2225 -291 2763
rect -17 2225 17 2763
rect 291 2225 325 2763
rect 599 2225 633 2763
rect -479 1826 -445 1860
rect -171 1826 -137 1860
rect 137 1826 171 1860
rect 445 1826 479 1860
rect -633 960 -599 1498
rect -325 960 -291 1498
rect -17 960 17 1498
rect 291 960 325 1498
rect 599 960 633 1498
rect -479 561 -445 595
rect -171 561 -137 595
rect 137 561 171 595
rect 445 561 479 595
rect -633 -305 -599 233
rect -325 -305 -291 233
rect -17 -305 17 233
rect 291 -305 325 233
rect 599 -305 633 233
rect -479 -704 -445 -670
rect -171 -704 -137 -670
rect 137 -704 171 -670
rect 445 -704 479 -670
rect -633 -1570 -599 -1032
rect -325 -1570 -291 -1032
rect -17 -1570 17 -1032
rect 291 -1570 325 -1032
rect 599 -1570 633 -1032
rect -479 -1969 -445 -1935
rect -171 -1969 -137 -1935
rect 137 -1969 171 -1935
rect 445 -1969 479 -1935
rect -633 -2835 -599 -2297
rect -325 -2835 -291 -2297
rect -17 -2835 17 -2297
rect 291 -2835 325 -2297
rect 599 -2835 633 -2297
<< metal1 >>
rect -491 3125 -433 3131
rect -491 3091 -479 3125
rect -445 3091 -433 3125
rect -491 3085 -433 3091
rect -183 3125 -125 3131
rect -183 3091 -171 3125
rect -137 3091 -125 3125
rect -183 3085 -125 3091
rect 125 3125 183 3131
rect 125 3091 137 3125
rect 171 3091 183 3125
rect 125 3085 183 3091
rect 433 3125 491 3131
rect 433 3091 445 3125
rect 479 3091 491 3125
rect 433 3085 491 3091
rect -639 2763 -593 2775
rect -639 2225 -633 2763
rect -599 2225 -593 2763
rect -639 2213 -593 2225
rect -331 2763 -285 2775
rect -331 2225 -325 2763
rect -291 2225 -285 2763
rect -331 2213 -285 2225
rect -23 2763 23 2775
rect -23 2225 -17 2763
rect 17 2225 23 2763
rect -23 2213 23 2225
rect 285 2763 331 2775
rect 285 2225 291 2763
rect 325 2225 331 2763
rect 285 2213 331 2225
rect 593 2763 639 2775
rect 593 2225 599 2763
rect 633 2225 639 2763
rect 593 2213 639 2225
rect -491 1860 -433 1866
rect -491 1826 -479 1860
rect -445 1826 -433 1860
rect -491 1820 -433 1826
rect -183 1860 -125 1866
rect -183 1826 -171 1860
rect -137 1826 -125 1860
rect -183 1820 -125 1826
rect 125 1860 183 1866
rect 125 1826 137 1860
rect 171 1826 183 1860
rect 125 1820 183 1826
rect 433 1860 491 1866
rect 433 1826 445 1860
rect 479 1826 491 1860
rect 433 1820 491 1826
rect -639 1498 -593 1510
rect -639 960 -633 1498
rect -599 960 -593 1498
rect -639 948 -593 960
rect -331 1498 -285 1510
rect -331 960 -325 1498
rect -291 960 -285 1498
rect -331 948 -285 960
rect -23 1498 23 1510
rect -23 960 -17 1498
rect 17 960 23 1498
rect -23 948 23 960
rect 285 1498 331 1510
rect 285 960 291 1498
rect 325 960 331 1498
rect 285 948 331 960
rect 593 1498 639 1510
rect 593 960 599 1498
rect 633 960 639 1498
rect 593 948 639 960
rect -491 595 -433 601
rect -491 561 -479 595
rect -445 561 -433 595
rect -491 555 -433 561
rect -183 595 -125 601
rect -183 561 -171 595
rect -137 561 -125 595
rect -183 555 -125 561
rect 125 595 183 601
rect 125 561 137 595
rect 171 561 183 595
rect 125 555 183 561
rect 433 595 491 601
rect 433 561 445 595
rect 479 561 491 595
rect 433 555 491 561
rect -639 233 -593 245
rect -639 -305 -633 233
rect -599 -305 -593 233
rect -639 -317 -593 -305
rect -331 233 -285 245
rect -331 -305 -325 233
rect -291 -305 -285 233
rect -331 -317 -285 -305
rect -23 233 23 245
rect -23 -305 -17 233
rect 17 -305 23 233
rect -23 -317 23 -305
rect 285 233 331 245
rect 285 -305 291 233
rect 325 -305 331 233
rect 285 -317 331 -305
rect 593 233 639 245
rect 593 -305 599 233
rect 633 -305 639 233
rect 593 -317 639 -305
rect -491 -670 -433 -664
rect -491 -704 -479 -670
rect -445 -704 -433 -670
rect -491 -710 -433 -704
rect -183 -670 -125 -664
rect -183 -704 -171 -670
rect -137 -704 -125 -670
rect -183 -710 -125 -704
rect 125 -670 183 -664
rect 125 -704 137 -670
rect 171 -704 183 -670
rect 125 -710 183 -704
rect 433 -670 491 -664
rect 433 -704 445 -670
rect 479 -704 491 -670
rect 433 -710 491 -704
rect -639 -1032 -593 -1020
rect -639 -1570 -633 -1032
rect -599 -1570 -593 -1032
rect -639 -1582 -593 -1570
rect -331 -1032 -285 -1020
rect -331 -1570 -325 -1032
rect -291 -1570 -285 -1032
rect -331 -1582 -285 -1570
rect -23 -1032 23 -1020
rect -23 -1570 -17 -1032
rect 17 -1570 23 -1032
rect -23 -1582 23 -1570
rect 285 -1032 331 -1020
rect 285 -1570 291 -1032
rect 325 -1570 331 -1032
rect 285 -1582 331 -1570
rect 593 -1032 639 -1020
rect 593 -1570 599 -1032
rect 633 -1570 639 -1032
rect 593 -1582 639 -1570
rect -491 -1935 -433 -1929
rect -491 -1969 -479 -1935
rect -445 -1969 -433 -1935
rect -491 -1975 -433 -1969
rect -183 -1935 -125 -1929
rect -183 -1969 -171 -1935
rect -137 -1969 -125 -1935
rect -183 -1975 -125 -1969
rect 125 -1935 183 -1929
rect 125 -1969 137 -1935
rect 171 -1969 183 -1935
rect 125 -1975 183 -1969
rect 433 -1935 491 -1929
rect 433 -1969 445 -1935
rect 479 -1969 491 -1935
rect 433 -1975 491 -1969
rect -639 -2297 -593 -2285
rect -639 -2835 -633 -2297
rect -599 -2835 -593 -2297
rect -639 -2847 -593 -2835
rect -331 -2297 -285 -2285
rect -331 -2835 -325 -2297
rect -291 -2835 -285 -2297
rect -331 -2847 -285 -2835
rect -23 -2297 23 -2285
rect -23 -2835 -17 -2297
rect 17 -2835 23 -2297
rect -23 -2847 23 -2835
rect 285 -2297 331 -2285
rect 285 -2835 291 -2297
rect 325 -2835 331 -2297
rect 285 -2847 331 -2835
rect 593 -2297 639 -2285
rect 593 -2835 599 -2297
rect 633 -2835 639 -2297
rect 593 -2847 639 -2835
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 5.5 l 1.25 m 5 nf 4 diffcov 50 polycov 20 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 class mosfet compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 50 viadrn 50 viagate 10 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1770979109
<< nwell >>
rect -423 -300 423 300
<< pmos >>
rect -329 -200 -29 200
rect 29 -200 329 200
<< pdiff >>
rect -387 188 -329 200
rect -387 -188 -375 188
rect -341 -188 -329 188
rect -387 -200 -329 -188
rect -29 188 29 200
rect -29 -188 -17 188
rect 17 -188 29 188
rect -29 -200 29 -188
rect 329 188 387 200
rect 329 -188 341 188
rect 375 -188 387 188
rect 329 -200 387 -188
<< pdiffc >>
rect -375 -188 -341 188
rect -17 -188 17 188
rect 341 -188 375 188
<< poly >>
rect -262 281 -96 297
rect -262 264 -246 281
rect -329 247 -246 264
rect -112 264 -96 281
rect 96 281 262 297
rect 96 264 112 281
rect -112 247 -29 264
rect -329 200 -29 247
rect 29 247 112 264
rect 246 264 262 281
rect 246 247 329 264
rect 29 200 329 247
rect -329 -247 -29 -200
rect -329 -264 -246 -247
rect -262 -281 -246 -264
rect -112 -264 -29 -247
rect 29 -247 329 -200
rect 29 -264 112 -247
rect -112 -281 -96 -264
rect -262 -297 -96 -281
rect 96 -281 112 -264
rect 246 -264 329 -247
rect 246 -281 262 -264
rect 96 -297 262 -281
<< polycont >>
rect -246 247 -112 281
rect 112 247 246 281
rect -246 -281 -112 -247
rect 112 -281 246 -247
<< locali >>
rect -262 247 -246 281
rect -112 247 -96 281
rect 96 247 112 281
rect 246 247 262 281
rect -375 188 -341 204
rect -375 -204 -341 -188
rect -17 188 17 204
rect -17 -204 17 -188
rect 341 188 375 204
rect 341 -204 375 -188
rect -262 -281 -246 -247
rect -112 -281 -96 -247
rect 96 -281 112 -247
rect 246 -281 262 -247
<< viali >>
rect -246 247 -112 281
rect 112 247 246 281
rect -375 -188 -341 188
rect -17 -188 17 188
rect 341 -188 375 188
rect -246 -281 -112 -247
rect 112 -281 246 -247
<< metal1 >>
rect -258 281 -100 287
rect -258 247 -246 281
rect -112 247 -100 281
rect -258 241 -100 247
rect 100 281 258 287
rect 100 247 112 281
rect 246 247 258 281
rect 100 241 258 247
rect -381 188 -335 200
rect -381 -188 -375 188
rect -341 -188 -335 188
rect -381 -200 -335 -188
rect -23 188 23 200
rect -23 -188 -17 188
rect 17 -188 23 188
rect -23 -200 23 -188
rect 335 188 381 200
rect 335 -188 341 188
rect 375 -188 381 188
rect 335 -200 381 -188
rect -258 -247 -100 -241
rect -258 -281 -246 -247
rect -112 -281 -100 -247
rect -258 -287 -100 -281
rect 100 -247 258 -241
rect 100 -281 112 -247
rect 246 -281 258 -247
rect 100 -287 258 -281
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 2.0 l 1.5 m 1 nf 2 diffcov 100 polycov 50 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 class mosfet compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 50 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

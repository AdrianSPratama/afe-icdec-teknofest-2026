magic
tech sky130A
magscale 1 2
timestamp 1771413069
<< error_p >>
rect -681 1915 681 2166
rect -681 650 681 901
rect -681 -615 681 -364
rect -681 -1880 681 -1629
<< nwell >>
rect -681 1915 681 3177
rect -681 650 681 1912
rect -681 -615 681 647
rect -681 -1880 681 -618
rect -681 -3145 681 -1883
<< pmos >>
rect -587 2015 -337 3115
rect -279 2015 -29 3115
rect 29 2015 279 3115
rect 337 2015 587 3115
rect -587 750 -337 1850
rect -279 750 -29 1850
rect 29 750 279 1850
rect 337 750 587 1850
rect -587 -515 -337 585
rect -279 -515 -29 585
rect 29 -515 279 585
rect 337 -515 587 585
rect -587 -1780 -337 -680
rect -279 -1780 -29 -680
rect 29 -1780 279 -680
rect 337 -1780 587 -680
rect -587 -3045 -337 -1945
rect -279 -3045 -29 -1945
rect 29 -3045 279 -1945
rect 337 -3045 587 -1945
<< pdiff >>
rect -645 3103 -587 3115
rect -645 2027 -633 3103
rect -599 2027 -587 3103
rect -645 2015 -587 2027
rect -337 3103 -279 3115
rect -337 2027 -325 3103
rect -291 2027 -279 3103
rect -337 2015 -279 2027
rect -29 3103 29 3115
rect -29 2027 -17 3103
rect 17 2027 29 3103
rect -29 2015 29 2027
rect 279 3103 337 3115
rect 279 2027 291 3103
rect 325 2027 337 3103
rect 279 2015 337 2027
rect 587 3103 645 3115
rect 587 2027 599 3103
rect 633 2027 645 3103
rect 587 2015 645 2027
rect -645 1838 -587 1850
rect -645 762 -633 1838
rect -599 762 -587 1838
rect -645 750 -587 762
rect -337 1838 -279 1850
rect -337 762 -325 1838
rect -291 762 -279 1838
rect -337 750 -279 762
rect -29 1838 29 1850
rect -29 762 -17 1838
rect 17 762 29 1838
rect -29 750 29 762
rect 279 1838 337 1850
rect 279 762 291 1838
rect 325 762 337 1838
rect 279 750 337 762
rect 587 1838 645 1850
rect 587 762 599 1838
rect 633 762 645 1838
rect 587 750 645 762
rect -645 573 -587 585
rect -645 -503 -633 573
rect -599 -503 -587 573
rect -645 -515 -587 -503
rect -337 573 -279 585
rect -337 -503 -325 573
rect -291 -503 -279 573
rect -337 -515 -279 -503
rect -29 573 29 585
rect -29 -503 -17 573
rect 17 -503 29 573
rect -29 -515 29 -503
rect 279 573 337 585
rect 279 -503 291 573
rect 325 -503 337 573
rect 279 -515 337 -503
rect 587 573 645 585
rect 587 -503 599 573
rect 633 -503 645 573
rect 587 -515 645 -503
rect -645 -692 -587 -680
rect -645 -1768 -633 -692
rect -599 -1768 -587 -692
rect -645 -1780 -587 -1768
rect -337 -692 -279 -680
rect -337 -1768 -325 -692
rect -291 -1768 -279 -692
rect -337 -1780 -279 -1768
rect -29 -692 29 -680
rect -29 -1768 -17 -692
rect 17 -1768 29 -692
rect -29 -1780 29 -1768
rect 279 -692 337 -680
rect 279 -1768 291 -692
rect 325 -1768 337 -692
rect 279 -1780 337 -1768
rect 587 -692 645 -680
rect 587 -1768 599 -692
rect 633 -1768 645 -692
rect 587 -1780 645 -1768
rect -645 -1957 -587 -1945
rect -645 -3033 -633 -1957
rect -599 -3033 -587 -1957
rect -645 -3045 -587 -3033
rect -337 -1957 -279 -1945
rect -337 -3033 -325 -1957
rect -291 -3033 -279 -1957
rect -337 -3045 -279 -3033
rect -29 -1957 29 -1945
rect -29 -3033 -17 -1957
rect 17 -3033 29 -1957
rect -29 -3045 29 -3033
rect 279 -1957 337 -1945
rect 279 -3033 291 -1957
rect 325 -3033 337 -1957
rect 279 -3045 337 -3033
rect 587 -1957 645 -1945
rect 587 -3033 599 -1957
rect 633 -3033 645 -1957
rect 587 -3045 645 -3033
<< pdiffc >>
rect -633 2027 -599 3103
rect -325 2027 -291 3103
rect -17 2027 17 3103
rect 291 2027 325 3103
rect 599 2027 633 3103
rect -633 762 -599 1838
rect -325 762 -291 1838
rect -17 762 17 1838
rect 291 762 325 1838
rect 599 762 633 1838
rect -633 -503 -599 573
rect -325 -503 -291 573
rect -17 -503 17 573
rect 291 -503 325 573
rect 599 -503 633 573
rect -633 -1768 -599 -692
rect -325 -1768 -291 -692
rect -17 -1768 17 -692
rect 291 -1768 325 -692
rect 599 -1768 633 -692
rect -633 -3033 -599 -1957
rect -325 -3033 -291 -1957
rect -17 -3033 17 -1957
rect 291 -3033 325 -1957
rect 599 -3033 633 -1957
<< poly >>
rect -587 3115 -337 3141
rect -279 3115 -29 3141
rect 29 3115 279 3141
rect 337 3115 587 3141
rect -587 1968 -337 2015
rect -587 1934 -571 1968
rect -353 1934 -337 1968
rect -587 1918 -337 1934
rect -279 1968 -29 2015
rect -279 1934 -263 1968
rect -45 1934 -29 1968
rect -279 1918 -29 1934
rect 29 1968 279 2015
rect 29 1934 45 1968
rect 263 1934 279 1968
rect 29 1918 279 1934
rect 337 1968 587 2015
rect 337 1934 353 1968
rect 571 1934 587 1968
rect 337 1918 587 1934
rect -587 1850 -337 1876
rect -279 1850 -29 1876
rect 29 1850 279 1876
rect 337 1850 587 1876
rect -587 703 -337 750
rect -587 669 -571 703
rect -353 669 -337 703
rect -587 653 -337 669
rect -279 703 -29 750
rect -279 669 -263 703
rect -45 669 -29 703
rect -279 653 -29 669
rect 29 703 279 750
rect 29 669 45 703
rect 263 669 279 703
rect 29 653 279 669
rect 337 703 587 750
rect 337 669 353 703
rect 571 669 587 703
rect 337 653 587 669
rect -587 585 -337 611
rect -279 585 -29 611
rect 29 585 279 611
rect 337 585 587 611
rect -587 -562 -337 -515
rect -587 -596 -571 -562
rect -353 -596 -337 -562
rect -587 -612 -337 -596
rect -279 -562 -29 -515
rect -279 -596 -263 -562
rect -45 -596 -29 -562
rect -279 -612 -29 -596
rect 29 -562 279 -515
rect 29 -596 45 -562
rect 263 -596 279 -562
rect 29 -612 279 -596
rect 337 -562 587 -515
rect 337 -596 353 -562
rect 571 -596 587 -562
rect 337 -612 587 -596
rect -587 -680 -337 -654
rect -279 -680 -29 -654
rect 29 -680 279 -654
rect 337 -680 587 -654
rect -587 -1827 -337 -1780
rect -587 -1861 -571 -1827
rect -353 -1861 -337 -1827
rect -587 -1877 -337 -1861
rect -279 -1827 -29 -1780
rect -279 -1861 -263 -1827
rect -45 -1861 -29 -1827
rect -279 -1877 -29 -1861
rect 29 -1827 279 -1780
rect 29 -1861 45 -1827
rect 263 -1861 279 -1827
rect 29 -1877 279 -1861
rect 337 -1827 587 -1780
rect 337 -1861 353 -1827
rect 571 -1861 587 -1827
rect 337 -1877 587 -1861
rect -587 -1945 -337 -1919
rect -279 -1945 -29 -1919
rect 29 -1945 279 -1919
rect 337 -1945 587 -1919
rect -587 -3092 -337 -3045
rect -587 -3126 -571 -3092
rect -353 -3126 -337 -3092
rect -587 -3142 -337 -3126
rect -279 -3092 -29 -3045
rect -279 -3126 -263 -3092
rect -45 -3126 -29 -3092
rect -279 -3142 -29 -3126
rect 29 -3092 279 -3045
rect 29 -3126 45 -3092
rect 263 -3126 279 -3092
rect 29 -3142 279 -3126
rect 337 -3092 587 -3045
rect 337 -3126 353 -3092
rect 571 -3126 587 -3092
rect 337 -3142 587 -3126
<< polycont >>
rect -571 1934 -353 1968
rect -263 1934 -45 1968
rect 45 1934 263 1968
rect 353 1934 571 1968
rect -571 669 -353 703
rect -263 669 -45 703
rect 45 669 263 703
rect 353 669 571 703
rect -571 -596 -353 -562
rect -263 -596 -45 -562
rect 45 -596 263 -562
rect 353 -596 571 -562
rect -571 -1861 -353 -1827
rect -263 -1861 -45 -1827
rect 45 -1861 263 -1827
rect 353 -1861 571 -1827
rect -571 -3126 -353 -3092
rect -263 -3126 -45 -3092
rect 45 -3126 263 -3092
rect 353 -3126 571 -3092
<< locali >>
rect -633 3103 -599 3119
rect -633 2011 -599 2027
rect -325 3103 -291 3119
rect -325 2011 -291 2027
rect -17 3103 17 3119
rect -17 2011 17 2027
rect 291 3103 325 3119
rect 291 2011 325 2027
rect 599 3103 633 3119
rect 599 2011 633 2027
rect -587 1934 -571 1968
rect -353 1934 -337 1968
rect -279 1934 -263 1968
rect -45 1934 -29 1968
rect 29 1934 45 1968
rect 263 1934 279 1968
rect 337 1934 353 1968
rect 571 1934 587 1968
rect -633 1838 -599 1854
rect -633 746 -599 762
rect -325 1838 -291 1854
rect -325 746 -291 762
rect -17 1838 17 1854
rect -17 746 17 762
rect 291 1838 325 1854
rect 291 746 325 762
rect 599 1838 633 1854
rect 599 746 633 762
rect -587 669 -571 703
rect -353 669 -337 703
rect -279 669 -263 703
rect -45 669 -29 703
rect 29 669 45 703
rect 263 669 279 703
rect 337 669 353 703
rect 571 669 587 703
rect -633 573 -599 589
rect -633 -519 -599 -503
rect -325 573 -291 589
rect -325 -519 -291 -503
rect -17 573 17 589
rect -17 -519 17 -503
rect 291 573 325 589
rect 291 -519 325 -503
rect 599 573 633 589
rect 599 -519 633 -503
rect -587 -596 -571 -562
rect -353 -596 -337 -562
rect -279 -596 -263 -562
rect -45 -596 -29 -562
rect 29 -596 45 -562
rect 263 -596 279 -562
rect 337 -596 353 -562
rect 571 -596 587 -562
rect -633 -692 -599 -676
rect -633 -1784 -599 -1768
rect -325 -692 -291 -676
rect -325 -1784 -291 -1768
rect -17 -692 17 -676
rect -17 -1784 17 -1768
rect 291 -692 325 -676
rect 291 -1784 325 -1768
rect 599 -692 633 -676
rect 599 -1784 633 -1768
rect -587 -1861 -571 -1827
rect -353 -1861 -337 -1827
rect -279 -1861 -263 -1827
rect -45 -1861 -29 -1827
rect 29 -1861 45 -1827
rect 263 -1861 279 -1827
rect 337 -1861 353 -1827
rect 571 -1861 587 -1827
rect -633 -1957 -599 -1941
rect -633 -3049 -599 -3033
rect -325 -1957 -291 -1941
rect -325 -3049 -291 -3033
rect -17 -1957 17 -1941
rect -17 -3049 17 -3033
rect 291 -1957 325 -1941
rect 291 -3049 325 -3033
rect 599 -1957 633 -1941
rect 599 -3049 633 -3033
rect -587 -3126 -571 -3092
rect -353 -3126 -337 -3092
rect -279 -3126 -263 -3092
rect -45 -3126 -29 -3092
rect 29 -3126 45 -3092
rect 263 -3126 279 -3092
rect 337 -3126 353 -3092
rect 571 -3126 587 -3092
<< viali >>
rect -633 2027 -599 3103
rect -325 2027 -291 3103
rect -17 2027 17 3103
rect 291 2027 325 3103
rect 599 2027 633 3103
rect -571 1934 -353 1968
rect -263 1934 -45 1968
rect 45 1934 263 1968
rect 353 1934 571 1968
rect -633 762 -599 1838
rect -325 762 -291 1838
rect -17 762 17 1838
rect 291 762 325 1838
rect 599 762 633 1838
rect -571 669 -353 703
rect -263 669 -45 703
rect 45 669 263 703
rect 353 669 571 703
rect -633 -503 -599 573
rect -325 -503 -291 573
rect -17 -503 17 573
rect 291 -503 325 573
rect 599 -503 633 573
rect -571 -596 -353 -562
rect -263 -596 -45 -562
rect 45 -596 263 -562
rect 353 -596 571 -562
rect -633 -1768 -599 -692
rect -325 -1768 -291 -692
rect -17 -1768 17 -692
rect 291 -1768 325 -692
rect 599 -1768 633 -692
rect -571 -1861 -353 -1827
rect -263 -1861 -45 -1827
rect 45 -1861 263 -1827
rect 353 -1861 571 -1827
rect -633 -3033 -599 -1957
rect -325 -3033 -291 -1957
rect -17 -3033 17 -1957
rect 291 -3033 325 -1957
rect 599 -3033 633 -1957
rect -571 -3126 -353 -3092
rect -263 -3126 -45 -3092
rect 45 -3126 263 -3092
rect 353 -3126 571 -3092
<< metal1 >>
rect -639 3103 -593 3115
rect -639 2027 -633 3103
rect -599 2027 -593 3103
rect -639 2015 -593 2027
rect -331 3103 -285 3115
rect -331 2027 -325 3103
rect -291 2027 -285 3103
rect -331 2015 -285 2027
rect -23 3103 23 3115
rect -23 2027 -17 3103
rect 17 2027 23 3103
rect -23 2015 23 2027
rect 285 3103 331 3115
rect 285 2027 291 3103
rect 325 2027 331 3103
rect 285 2015 331 2027
rect 593 3103 639 3115
rect 593 2027 599 3103
rect 633 2027 639 3103
rect 593 2015 639 2027
rect -583 1968 -341 1974
rect -583 1934 -571 1968
rect -353 1934 -341 1968
rect -583 1928 -341 1934
rect -275 1968 -33 1974
rect -275 1934 -263 1968
rect -45 1934 -33 1968
rect -275 1928 -33 1934
rect 33 1968 275 1974
rect 33 1934 45 1968
rect 263 1934 275 1968
rect 33 1928 275 1934
rect 341 1968 583 1974
rect 341 1934 353 1968
rect 571 1934 583 1968
rect 341 1928 583 1934
rect -639 1838 -593 1850
rect -639 762 -633 1838
rect -599 762 -593 1838
rect -639 750 -593 762
rect -331 1838 -285 1850
rect -331 762 -325 1838
rect -291 762 -285 1838
rect -331 750 -285 762
rect -23 1838 23 1850
rect -23 762 -17 1838
rect 17 762 23 1838
rect -23 750 23 762
rect 285 1838 331 1850
rect 285 762 291 1838
rect 325 762 331 1838
rect 285 750 331 762
rect 593 1838 639 1850
rect 593 762 599 1838
rect 633 762 639 1838
rect 593 750 639 762
rect -583 703 -341 709
rect -583 669 -571 703
rect -353 669 -341 703
rect -583 663 -341 669
rect -275 703 -33 709
rect -275 669 -263 703
rect -45 669 -33 703
rect -275 663 -33 669
rect 33 703 275 709
rect 33 669 45 703
rect 263 669 275 703
rect 33 663 275 669
rect 341 703 583 709
rect 341 669 353 703
rect 571 669 583 703
rect 341 663 583 669
rect -639 573 -593 585
rect -639 -503 -633 573
rect -599 -503 -593 573
rect -639 -515 -593 -503
rect -331 573 -285 585
rect -331 -503 -325 573
rect -291 -503 -285 573
rect -331 -515 -285 -503
rect -23 573 23 585
rect -23 -503 -17 573
rect 17 -503 23 573
rect -23 -515 23 -503
rect 285 573 331 585
rect 285 -503 291 573
rect 325 -503 331 573
rect 285 -515 331 -503
rect 593 573 639 585
rect 593 -503 599 573
rect 633 -503 639 573
rect 593 -515 639 -503
rect -583 -562 -341 -556
rect -583 -596 -571 -562
rect -353 -596 -341 -562
rect -583 -602 -341 -596
rect -275 -562 -33 -556
rect -275 -596 -263 -562
rect -45 -596 -33 -562
rect -275 -602 -33 -596
rect 33 -562 275 -556
rect 33 -596 45 -562
rect 263 -596 275 -562
rect 33 -602 275 -596
rect 341 -562 583 -556
rect 341 -596 353 -562
rect 571 -596 583 -562
rect 341 -602 583 -596
rect -639 -692 -593 -680
rect -639 -1768 -633 -692
rect -599 -1768 -593 -692
rect -639 -1780 -593 -1768
rect -331 -692 -285 -680
rect -331 -1768 -325 -692
rect -291 -1768 -285 -692
rect -331 -1780 -285 -1768
rect -23 -692 23 -680
rect -23 -1768 -17 -692
rect 17 -1768 23 -692
rect -23 -1780 23 -1768
rect 285 -692 331 -680
rect 285 -1768 291 -692
rect 325 -1768 331 -692
rect 285 -1780 331 -1768
rect 593 -692 639 -680
rect 593 -1768 599 -692
rect 633 -1768 639 -692
rect 593 -1780 639 -1768
rect -583 -1827 -341 -1821
rect -583 -1861 -571 -1827
rect -353 -1861 -341 -1827
rect -583 -1867 -341 -1861
rect -275 -1827 -33 -1821
rect -275 -1861 -263 -1827
rect -45 -1861 -33 -1827
rect -275 -1867 -33 -1861
rect 33 -1827 275 -1821
rect 33 -1861 45 -1827
rect 263 -1861 275 -1827
rect 33 -1867 275 -1861
rect 341 -1827 583 -1821
rect 341 -1861 353 -1827
rect 571 -1861 583 -1827
rect 341 -1867 583 -1861
rect -639 -1957 -593 -1945
rect -639 -3033 -633 -1957
rect -599 -3033 -593 -1957
rect -639 -3045 -593 -3033
rect -331 -1957 -285 -1945
rect -331 -3033 -325 -1957
rect -291 -3033 -285 -1957
rect -331 -3045 -285 -3033
rect -23 -1957 23 -1945
rect -23 -3033 -17 -1957
rect 17 -3033 23 -1957
rect -23 -3045 23 -3033
rect 285 -1957 331 -1945
rect 285 -3033 291 -1957
rect 325 -3033 331 -1957
rect 285 -3045 331 -3033
rect 593 -1957 639 -1945
rect 593 -3033 599 -1957
rect 633 -3033 639 -1957
rect 593 -3045 639 -3033
rect -583 -3092 -341 -3086
rect -583 -3126 -571 -3092
rect -353 -3126 -341 -3092
rect -583 -3132 -341 -3126
rect -275 -3092 -33 -3086
rect -275 -3126 -263 -3092
rect -45 -3126 -33 -3092
rect -275 -3132 -33 -3126
rect 33 -3092 275 -3086
rect 33 -3126 45 -3092
rect 263 -3126 275 -3092
rect 33 -3132 275 -3126
rect 341 -3092 583 -3086
rect 341 -3126 353 -3092
rect 571 -3126 583 -3092
rect 341 -3132 583 -3126
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 5.5 l 1.25 m 5 nf 4 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 class mosfet compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

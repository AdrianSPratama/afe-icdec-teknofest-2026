magic
tech sky130A
magscale 1 2
timestamp 1771413069
<< nwell >>
rect -681 -334 681 368
<< pmos >>
rect -587 -234 -337 306
rect -279 -234 -29 306
rect 29 -234 279 306
rect 337 -234 587 306
<< pdiff >>
rect -645 294 -587 306
rect -645 -222 -633 294
rect -599 -222 -587 294
rect -645 -234 -587 -222
rect -337 294 -279 306
rect -337 -222 -325 294
rect -291 -222 -279 294
rect -337 -234 -279 -222
rect -29 294 29 306
rect -29 -222 -17 294
rect 17 -222 29 294
rect -29 -234 29 -222
rect 279 294 337 306
rect 279 -222 291 294
rect 325 -222 337 294
rect 279 -234 337 -222
rect 587 294 645 306
rect 587 -222 599 294
rect 633 -222 645 294
rect 587 -234 645 -222
<< pdiffc >>
rect -633 -222 -599 294
rect -325 -222 -291 294
rect -17 -222 17 294
rect 291 -222 325 294
rect 599 -222 633 294
<< poly >>
rect -587 306 -337 332
rect -279 306 -29 332
rect 29 306 279 332
rect 337 306 587 332
rect -587 -281 -337 -234
rect -587 -315 -571 -281
rect -353 -315 -337 -281
rect -587 -331 -337 -315
rect -279 -281 -29 -234
rect -279 -315 -263 -281
rect -45 -315 -29 -281
rect -279 -331 -29 -315
rect 29 -281 279 -234
rect 29 -315 45 -281
rect 263 -315 279 -281
rect 29 -331 279 -315
rect 337 -281 587 -234
rect 337 -315 353 -281
rect 571 -315 587 -281
rect 337 -331 587 -315
<< polycont >>
rect -571 -315 -353 -281
rect -263 -315 -45 -281
rect 45 -315 263 -281
rect 353 -315 571 -281
<< locali >>
rect -633 294 -599 310
rect -633 -238 -599 -222
rect -325 294 -291 310
rect -325 -238 -291 -222
rect -17 294 17 310
rect -17 -238 17 -222
rect 291 294 325 310
rect 291 -238 325 -222
rect 599 294 633 310
rect 599 -238 633 -222
rect -587 -315 -571 -281
rect -353 -315 -337 -281
rect -279 -315 -263 -281
rect -45 -315 -29 -281
rect 29 -315 45 -281
rect 263 -315 279 -281
rect 337 -315 353 -281
rect 571 -315 587 -281
<< viali >>
rect -633 -222 -599 294
rect -325 -222 -291 294
rect -17 -222 17 294
rect 291 -222 325 294
rect 599 -222 633 294
rect -571 -315 -353 -281
rect -263 -315 -45 -281
rect 45 -315 263 -281
rect 353 -315 571 -281
<< metal1 >>
rect -639 294 -593 306
rect -639 -222 -633 294
rect -599 -222 -593 294
rect -639 -234 -593 -222
rect -331 294 -285 306
rect -331 -222 -325 294
rect -291 -222 -285 294
rect -331 -234 -285 -222
rect -23 294 23 306
rect -23 -222 -17 294
rect 17 -222 23 294
rect -23 -234 23 -222
rect 285 294 331 306
rect 285 -222 291 294
rect 325 -222 331 294
rect 285 -234 331 -222
rect 593 294 639 306
rect 593 -222 599 294
rect 633 -222 639 294
rect 593 -234 639 -222
rect -583 -281 -341 -275
rect -583 -315 -571 -281
rect -353 -315 -341 -281
rect -583 -321 -341 -315
rect -275 -281 -33 -275
rect -275 -315 -263 -281
rect -45 -315 -33 -281
rect -275 -321 -33 -315
rect 33 -281 275 -275
rect 33 -315 45 -281
rect 263 -315 275 -281
rect 33 -321 275 -315
rect 341 -281 583 -275
rect 341 -315 353 -281
rect 571 -315 583 -281
rect 341 -321 583 -315
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 2.7 l 1.25 m 1 nf 4 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 class mosfet compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
